-- ---------------------------------------------------------------------
-- @file : uCore.vhd
-- ---------------------------------------------------------------------
--
-- Last change: KS 04.03.2021 16:46:38
-- Project : microCore
-- Language : VHDL-2008
-- Last check in : $Rev: 664 $ $Date:: 2021-03-10 #$
-- @copyright (c): Klaus Schleisiek, All Rights Reserved.
--
-- Do not use this file except in compliance with the License.
-- You may obtain a copy of the License at
-- https://github.com/microCore-VHDL/microCore/tree/master/documents
-- Software distributed under the License is distributed on an "AS IS"
-- basis, WITHOUT WARRANTY OF ANY KIND, either express or implied.
-- See the License for the specific language governing rights and
-- limitations under the License.
--
-- @brief: The microCore processor kernel.
--
-- Version Author   Date       Changes
--   210     ks    8-Jun-2020  initial version
--   2300    ks    8-Mar-2021  compiler switch WITH_PROG_RW eliminated
--                             Conversion to NUMERIC_STD
-- ---------------------------------------------------------------------
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
USE work.functions_pkg.ALL;
USE work.architecture_pkg.ALL;

ENTITY microcore IS PORT (
   uBus        : IN    uBus_port;
   core        : OUT   core_signals;
   ext_memory  : OUT   datamem_port;
   ext_rdata   : IN    data_bus;
   dma         : IN    datamem_port;
   dma_rdata   : OUT   data_bus;
-- umbilical uart interface
   rxd         : IN    STD_LOGIC;
   break       : OUT   STD_LOGIC;
   txd         : OUT   STD_LOGIC
); END microcore;

ARCHITECTURE rtl OF microcore IS

ATTRIBUTE syn_keep  : BOOLEAN;
ATTRIBUTE init      : STRING;

ALIAS  reset     : STD_LOGIC IS uBus.reset;
ALIAS  clk       : STD_LOGIC IS uBus.clk;
ALIAS  clk_en    : STD_LOGIC IS uBus.clk_en;
ALIAS  delay     : STD_LOGIC IS uBus.delay;
ALIAS  pause     : STD_LOGIC IS uBus.pause;

SIGNAL cycle_ctr : NATURAL RANGE 0 TO cycles - 1;

COMPONENT microcontrol PORT (
   uBus        : IN  uBus_port;
   deb_reset   : IN  STD_LOGIC;    -- reset issued by debugger
   deb_pause   : IN  STD_LOGIC;    -- pause issued by debugger
   deb_penable : IN  STD_LOGIC;    -- program memory ready for write by debugger
   uCtrl       : OUT core_signals;
   progmem     : OUT progmem_port;
   prog_rdata  : IN  inst_bus;
   datamem		: OUT datamem_port;
   mem_rdata   : IN  data_bus      -- data memory read data
); END COMPONENT microcontrol;

SIGNAL uCtrl        : core_signals;
SIGNAL progmem      : progmem_port;
SIGNAL prog_rdata   : inst_bus;
SIGNAL datamem      : datamem_port;
SIGNAL memory       : datamem_port;
SIGNAL mem_rdata    : data_bus;

COMPONENT debugger PORT (
   uBus           : IN  uBus_port;
   deb_reset      : OUT STD_LOGIC;    -- reset generated by debugger
   deb_pause      : OUT STD_LOGIC;
   deb_prequest   : OUT STD_LOGIC;    -- request program memory write cycle
   deb_penable    : IN  STD_LOGIC;    -- execute program memory write
   deb_drequest   : OUT STD_LOGIC;    -- request data memory for a read/write cycle
   deb_denable    : IN  STD_LOGIC;    -- execute data memory read/write
   umbilical      : OUT progmem_port; -- interface to the program memory
   debugmem       : OUT datamem_port; -- interface to the data memory
   debugmem_rdata : IN  data_bus;
-- umbilical uart
   rxd            : IN  STD_LOGIC;
   break          : OUT STD_LOGIC;
   txd            : OUT STD_LOGIC
); END COMPONENT debugger;

SIGNAL umbilical     : progmem_port;
SIGNAL debugmem      : datamem_port;
SIGNAL deb_pause     : STD_LOGIC;
SIGNAL deb_reset     : STD_LOGIC;
SIGNAL deb_prequest  : STD_LOGIC;
SIGNAL deb_drequest  : STD_LOGIC;
SIGNAL deb_penable   : STD_LOGIC;
SIGNAL deb_denable   : STD_LOGIC;

SIGNAL warmboot      : STD_LOGIC := '0';
   ATTRIBUTE syn_keep OF warmboot : SIGNAL IS true;
   ATTRIBUTE init     OF warmboot : SIGNAL IS "0";

-- cold boot loader
COMPONENT boot_rom PORT (
   addr  : IN   boot_addr_bus;
   data  : OUT  inst_bus
); END COMPONENT boot_rom;

SIGNAL boot_addr   : boot_addr_bus;
SIGNAL boot_rdata  : inst_bus;

-- data memory
COMPONENT uDatacache PORT (
   clk          : IN  STD_LOGIC;
   enable       : IN  STD_LOGIC;
   write        : IN  STD_LOGIC;
   addr         : IN  dcache_addr;
   wdata        : IN  data_bus;
   rdata        : OUT data_bus;
   dma_enable   : IN  STD_LOGIC;
   dma_write    : IN  STD_LOGIC;
   dma_addr     : IN  dcache_addr;
   dma_wdata    : IN  data_bus;
   dma_rdata    : OUT data_bus
); END COMPONENT uDatacache;

SIGNAL dcache_en      : STD_LOGIC;
SIGNAL dcache_rdata   : data_bus;
SIGNAL ext_mem_en     : STD_LOGIC;
SIGNAL mem_addr       : data_addr;

-- program memory
COMPONENT uProgmem PORT (
   clk      : IN  STD_LOGIC;
   penable  : IN  STD_LOGIC;
   pwrite   : IN  STD_LOGIC;
   paddr    : IN  program_addr;
   pwdata   : IN  inst_bus;
   prdata   : OUT inst_bus
); END COMPONENT uProgmem;

SIGNAL pcache_rdata   : inst_bus;
SIGNAL pcache_wdata   : inst_bus;
SIGNAL pwrite         : STD_LOGIC;
SIGNAL paddr          : program_addr;

BEGIN

-- make sure reg_addr_width is large enough for all registers
ASSERT ((-1 * min_registers) < (2 ** reg_addr_width-1))
REPORT "reg_addr_width too small"
SEVERITY error;

-- ---------------------------------------------------------------------
-- sub-uCore cycle control
-- ---------------------------------------------------------------------

enable_proc: PROCESS (clk)
BEGIN
   IF  rising_edge(clk)  THEN
      IF  cycle_ctr = 0  THEN
         IF  delay = '0'  THEN
            cycle_ctr <= cycles - 1;
         END IF;
      ELSE
         cycle_ctr <= cycle_ctr - 1;
      END IF;
   END IF;
END PROCESS enable_proc;

-- ---------------------------------------------------------------------
-- internal data memory
-- ---------------------------------------------------------------------

memory <= debugmem WHEN  deb_denable = '1'  ELSE datamem;

with_ext_mem: IF  data_addr_width > cache_addr_width  GENERATE

   ext_mem_en <= '1' WHEN  uCtrl.ext_en = '1' OR
                           (deb_denable = '1' AND debugmem.addr(data_addr_width-1 DOWNTO cache_addr_width) /= 0)
                 ELSE '0';

END GENERATE with_ext_mem; no_ext_mem: IF  data_addr_width <= cache_addr_width  GENERATE

   ext_mem_en <= '0';

END GENERATE no_ext_mem;

ext_memory.enable <= ext_mem_en;
ext_memory.write  <= memory.write;
ext_memory.addr   <= memory.addr;
ext_memory.wdata  <= memory.wdata;

dcache_en <= clk_en AND NOT ext_mem_en AND memory.enable;

internal_data_mem: uDatacache PORT MAP (
   clk          => clk,
   enable       => dcache_en,
   write        => memory.write,
   addr         => memory.addr(cache_addr_width-1 DOWNTO 0),
   wdata        => memory.wdata,
   rdata        => dcache_rdata,
   dma_enable   => dma.enable,
   dma_write    => dma.write,
   dma_addr     => dma.addr(cache_addr_width-1 DOWNTO 0),
   dma_wdata    => dma.wdata,
   dma_rdata    => dma_rdata
);

-- pragma translate_off
memaddr_proc : PROCESS (clk)
BEGIN
   IF  rising_edge(clk)  THEN
      IF  dcache_en = '1'  THEN
         mem_addr <= memory.addr; -- state of the internal blockRAM address register for simulation
      END IF;
END IF;
END PROCESS memaddr_proc;
-- pragma translate_on

mem_rdata <= ext_rdata WHEN  ext_mem_en = '1'  ELSE  dcache_rdata;

-- ---------------------------------------------------------------------
-- internal program memory
-- ---------------------------------------------------------------------

paddr <= umbilical.addr  WHEN  deb_penable = '1'  ELSE  progmem.addr;

pwrite <= umbilical.write WHEN  deb_penable = '1'             ELSE
          progmem.write   WHEN  warmboot = '0' OR SIMULATION  ELSE '0'; -- only during boot phase

pcache_wdata <= umbilical.wdata  WHEN  deb_penable = '1'  ELSE  progmem.wdata;

internal_prog_mem: uProgmem PORT MAP (
   clk      => clk,
   penable  => clk_en,
   pwrite   => pwrite,
   paddr    => paddr,
   pwdata   => pcache_wdata,
   prdata   => pcache_rdata
);

prog_rdata <= pcache_rdata WHEN  warmboot = '1'  ELSE boot_rdata;

-- ---------------------------------------------------------------------
-- boot loader, reads from program memory after branch to zero (reboot)
-- ---------------------------------------------------------------------

cold_boot_proc: PROCESS (reset, clk)
BEGIN
   IF  reset = '1' AND async_reset  THEN
      IF  coldboot  THEN  warmboot <= '0';  END IF; -- go into boot loading on reset?
      boot_addr <= (OTHERS => '0');
   ELSIF  rising_edge(clk)  THEN
      IF  clk_en = '1' AND warmboot = '0'  THEN
         boot_addr <= progmem.addr(boot_addr_width-1 DOWNTO 0);
         IF  (prog_rdata = op_BRANCH AND progmem.addr = 0 AND progmem.write = '0') OR deb_penable = '1'  THEN
            warmboot <= '1';
         END IF;
      END IF;
      IF  reset = '1' AND NOT async_reset  THEN
         IF  coldboot  THEN  warmboot <= '0';  END IF; -- go into boot loading on reset?
         boot_addr <= (OTHERS => '0');
      END IF;
   END IF;
END PROCESS cold_boot_proc;

boot_loader: boot_rom PORT MAP(boot_addr, boot_rdata);

-- ---------------------------------------------------------------------
-- instruction execution engine
-- ---------------------------------------------------------------------

uCntrl: microcontrol PORT MAP (
   uBus        => uBus,
   deb_reset   => deb_reset,   -- reset issued by debugger
   deb_pause   => deb_pause,   -- pause issued by debugger
   deb_penable => deb_penable, -- program memory ready for write by debugger
   uCtrl       => uCtrl,
   progmem     => progmem,
   prog_rdata  => prog_rdata,
   datamem     => datamem,
   mem_rdata   => mem_rdata
);

core.clk_en    <= '1' WHEN  delay = '0' AND cycle_ctr = 0  ELSE '0';
core.reg_en    <= uCtrl.reg_en;
core.reg_addr  <= uCtrl.reg_addr;
core.ext_en    <= uCtrl.ext_en;
core.tick      <= uCtrl.tick;
core.chain     <= uCtrl.chain;
core.status    <= uCtrl.status;
core.dsp       <= uCtrl.dsp;
core.rsp       <= uCtrl.rsp;
core.int       <= uCtrl.int;
core.time      <= uCtrl.time;
core.debug     <= debugmem.wdata;

-- ---------------------------------------------------------------------
-- umbilical uart debug interface
-- ---------------------------------------------------------------------

deb_penable <= deb_prequest AND (NOT uCtrl.chain OR deb_reset);

deb_denable <= deb_drequest AND NOT (uCtrl.chain OR datamem.enable OR uCtrl.ext_en);

debug_unit: debugger PORT MAP (
   uBus           => uBus,
   deb_reset      => deb_reset,
   deb_pause      => deb_pause,
   deb_prequest   => deb_prequest,
   deb_penable    => deb_penable,
   deb_drequest   => deb_drequest,
   deb_denable    => deb_denable,
   umbilical      => umbilical,
   debugmem       => debugmem,
   debugmem_rdata => mem_rdata,
-- umbilical
   rxd            => rxd,
   break          => break,
   txd            => txd
);

END rtl;