-- ---------------------------------------------------------------------
-- @file : uDatacache_16b.vhd
-- ---------------------------------------------------------------------
--
-- Last change: KS 02.11.2022 23:17:05
-- @project: microCore
-- @language: VHDL-93
-- @copyright (c): Klaus Schleisiek, All Rights Reserved.
-- @contributors:
--
-- @license: Do not use this file except in compliance with the License.
-- You may obtain a copy of the Public License at
-- https://github.com/microCore-VHDL/microCore/tree/master/documents
-- Software distributed under the License is distributed on an "AS IS"
-- basis, WITHOUT WARRANTY OF ANY KIND, either express or implied.
-- See the License for the specific language governing rights and
-- limitations under the License.
--
-- @brief: Definition of the internal data memory.
-- Here fpga specific dual port memory IP for 16 bits has been included.
-- Parameters for 32 bits are:
-- CONSTANT data_width         : NATURAL := 32; -- data bus width
-- CONSTANT cache_size         : NATURAL := 16#C00#; -- data cache memory size
-- CONSTANT addr_rstack        : NATURAL := 16#800#; -- beginning of the return stack, must be a multiple of 2**rsp_width
--
-- Version Author   Date       Changes
--   210     ks    8-Jun-2020  initial version
--  2300     ks    8-Mar-2021  Conversion to NUMERIC_STD
--  2400     ks   03-Nov-2022  byte addressing using byte_addr_width > 0
-- ---------------------------------------------------------------------
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
USE work.functions_pkg.ALL;
USE work.architecture_pkg.ALL;

ENTITY uDatacache IS PORT (
   uBus        : IN  uBus_port;
   rdata       : OUT data_bus;
   dma_mem     : IN  datamem_port;
   dma_rdata   : OUT data_bus
); END uDatacache;

ARCHITECTURE rtl OF uDatacache IS

ALIAS clk            : STD_LOGIC IS uBus.clk;
ALIAS clk_en         : STD_LOGIC IS uBus.clk_en;
ALIAS mem_en         : STD_LOGIC IS uBus.mem_en;
ALIAS bytes          : byte_type IS uBus.bytes;
ALIAS write          : STD_LOGIC IS uBus.write;
ALIAS addr           : data_addr IS uBus.addr;
ALIAS wdata          : data_bus  IS uBus.wdata;
ALIAS dma_enable     : STD_LOGIC IS dma_mem.enable;
ALIAS dma_bytes      : byte_type IS dma_mem.bytes;
ALIAS dma_write      : STD_LOGIC IS dma_mem.write;
ALIAS dma_addr       : data_addr IS dma_mem.addr;
ALIAS dma_wdata      : data_bus  IS dma_mem.wdata;

SIGNAL enable        : STD_LOGIC;

SIGNAL bytes_en      : byte_addr;
SIGNAL mem_wdata     : data_bus;
SIGNAL mem_rdata     : data_bus;

SIGNAL dma_bytes_en  : byte_addr;
SIGNAL dma_mem_wdata : data_bus;
SIGNAL dma_mem_rdata : data_bus;

-- internal_datamem has been generated by IP-Express, Memory, EBR with the following parameters:
-- RAM_DP_TRUE, Depth 6144, Width 16, Normal, Big-Endian, ByteEn
COMPONENT byte_cache_16 PORT (
   ResetA    : IN  STD_LOGIC;
   ClockA    : IN  STD_LOGIC;
   ClockEnA  : IN  STD_LOGIC;
   WrA       : IN  STD_LOGIC;
   ByteEnA   : IN  STD_LOGIC_VECTOR(1 DOWNTO 0);
   AddressA  : IN  STD_LOGIC_VECTOR(12 DOWNTO 0);
   DataInA   : IN  STD_LOGIC_VECTOR(15 DOWNTO 0);
   QA        : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
-- dma port
   ResetB    : IN  STD_LOGIC;
   ClockB    : IN  STD_LOGIC;
   ClockEnB  : IN  STD_LOGIC;
   WrB       : IN  STD_LOGIC;
   ByteEnB   : IN  STD_LOGIC_VECTOR(1 DOWNTO 0);
   AddressB  : IN  STD_LOGIC_VECTOR(12 DOWNTO 0);
   DataInB   : IN  STD_LOGIC_VECTOR(15 DOWNTO 0);
   QB        : OUT STD_LOGIC_VECTOR(15 DOWNTO 0));
END COMPONENT byte_cache_16;

SIGNAL slv_mem_rdata  : STD_LOGIC_VECTOR(rdata'range);
SIGNAL slv_dma_rdata  : STD_LOGIC_VECTOR(dma_rdata'range);

BEGIN

enable <= clk_en AND mem_en;

byte_access_proc : PROCESS(uBus, mem_rdata, addr, dma_mem, dma_mem_rdata, dma_addr, bytes)
BEGIN

   mem_wdata <= wdata;
   rdata <= mem_rdata;
   bytes_en <= (OTHERS => '1');

   dma_mem_wdata <= dma_wdata;
   dma_rdata <= dma_mem_rdata;
   dma_bytes_en <= (OTHERS => '1');

-- 16 bit system
   IF  byte_addr_width = 1  THEN
      IF  bytes = 1  THEN        -- byte access
         mem_wdata <= wdata(7 DOWNTO 0) & wdata(7 DOWNTO  0);
         bytes_en <= "01";
         rdata <= resize(mem_rdata(07 DOWNTO 0), data_width);
         IF  addr(0) = '1'  THEN
            bytes_en <= "10";
            rdata <= resize(mem_rdata(15 DOWNTO 8), data_width);
         END IF;
         dma_mem_wdata <= dma_wdata(7 DOWNTO 0) & dma_wdata(7 DOWNTO  0);
         dma_bytes_en <= "01";
         dma_rdata <= resize(dma_mem_rdata(07 DOWNTO 0), data_width);
         IF  dma_addr(0) = '1'  THEN
            dma_bytes_en <= "10";
            dma_rdata <= resize(dma_mem_rdata(15 DOWNTO 8), data_width);
         END IF;
      END IF;
   END IF;

-- 32 bit system
   IF  byte_addr_width = 2  THEN
      IF  bytes = 1  THEN           -- byte access
         mem_wdata <= wdata(7 DOWNTO  0) & wdata(7 DOWNTO  0) & wdata(7 DOWNTO  0) & wdata(7 DOWNTO  0);
         CASE addr(1 DOWNTO 0) IS
         WHEN "00" => bytes_en <= "0001";
                      rdata <= resize(mem_rdata(07 DOWNTO 00), data_width);
         WHEN "01" => bytes_en <= "0010";
                      rdata <= resize(mem_rdata(15 DOWNTO 08), data_width);
         WHEN "10" => bytes_en <= "0100";
                      rdata <= resize(mem_rdata(23 DOWNTO 16), data_width);
         WHEN "11" => bytes_en <= "1000";
                      rdata <= resize(mem_rdata(31 DOWNTO 24), data_width);
         WHEN OTHERS => NULL;
         END CASE;
         dma_mem_wdata <= dma_wdata( 7 DOWNTO  0) & dma_wdata( 7 DOWNTO  0) & dma_wdata( 7 DOWNTO  0) & dma_wdata( 7 DOWNTO  0);
         CASE dma_addr(1 DOWNTO 0) IS
         WHEN "00" => dma_bytes_en <= "0001";
                      dma_rdata <= resize(dma_mem_rdata(07 DOWNTO 00), data_width);
         WHEN "01" => dma_bytes_en <= "0010";
                      dma_rdata <= resize(dma_mem_rdata(15 DOWNTO 08), data_width);
         WHEN "10" => dma_bytes_en <= "0100";
                      dma_rdata <= resize(dma_mem_rdata(23 DOWNTO 16), data_width);
         WHEN "11" => dma_bytes_en <= "1000";
                      dma_rdata <= resize(dma_mem_rdata(31 DOWNTO 24), data_width);
         WHEN OTHERS => NULL;
         END CASE;
      ELSIF  bytes = 2  THEN         -- word access
         mem_wdata <= wdata(15 DOWNTO 0) & wdata(15 DOWNTO  0);
         bytes_en <= "0011";
         rdata <= resize(mem_rdata(15 DOWNTO 0), data_width);
         IF  addr(1) = '1'  THEN
            bytes_en <= "1100";
            rdata <= resize(mem_rdata(31 DOWNTO 16), data_width);
         END IF;
         dma_mem_wdata <= dma_wdata(15 DOWNTO 0) & dma_wdata(15 DOWNTO  0);
         dma_bytes_en <= "0011";
         dma_rdata <= resize(dma_mem_rdata(15 DOWNTO 0), data_width);
         IF  dma_addr(1) = '1'  THEN
            dma_bytes_en <= "1100";
            dma_rdata <= resize(dma_mem_rdata(31 DOWNTO 16), data_width);
         END IF;
      END IF;
   END IF;

END PROCESS byte_access_proc;

make_sim_mem: IF  SIMULATION  GENERATE

   internal_data_mem: internal_dpbram
   GENERIC MAP (data_width, cache_size, byte_addr_width, "rw_check", DMEM_file)
   PORT MAP (
      clk     => clk,
      ena     => enable,
      wea     => write,
      bytea   => bytes_en,
      addra   => addr(cache_addr_width-1 DOWNTO byte_addr_width),
      dia     => mem_wdata,
      doa     => mem_rdata,
   -- dma port
      enb     => dma_enable,
      web     => dma_write,
      byteb   => dma_bytes_en,
      addrb   => dma_addr(cache_addr_width-1 DOWNTO byte_addr_width),
      dib     => dma_mem_wdata,
      dob     => dma_mem_rdata
   );

END GENERATE make_sim_mem; make_syn_mem: IF  NOT SIMULATION  GENERATE
-- instantiate FPGA specific IP for byte addressed memory here:

   instantiated_data_mem: byte_cache_16
   PORT MAP (
      ResetA    => '0',
      ClockA    => clk,
      ClockEnA  => enable,
      WrA       => write,
      ByteEnA   => std_logic_vector(bytes_en),
      AddressA  => std_logic_vector(addr(cache_addr_width-1 DOWNTO byte_addr_width)),
      DataInA   => std_logic_vector(mem_wdata),
      QA        => slv_mem_rdata,
-- dma port
      ResetB    => '0',
      ClockB    => clk,
      ClockEnB  => dma_enable,
      WrB       => dma_write,
      ByteEnB   => std_logic_vector(dma_bytes_en),
      AddressB  => std_logic_vector(dma_addr(cache_addr_width-1 DOWNTO byte_addr_width)),
      DataInB   => std_logic_vector(dma_mem_wdata),
      QB        => slv_dma_rdata
	);

   mem_rdata     <= unsigned(slv_mem_rdata);
   dma_mem_rdata <= unsigned(slv_dma_rdata);

END GENERATE make_syn_mem;

END rtl;

-- VHDL netlist generated by SCUBA Diamond (64-bit) 3.11.3.469
-- Module  Version: 7.5
--C:\lscc\diamond\3.11_x64\ispfpga\bin\nt64\scuba.exe -w -n byte_cache_16 -lang vhdl -synth synplify -bus_exp 7 -bb -arch mg5a00 -type bram -wp 11 -rp 1010
-- -data_width 16 -rdata_width 16 -num_rows 6144 -byte 8 -outdataB REGISTERED -writemodeA NORMAL -writemodeB NORMAL -resetmode SYNC -cascade -1

-- Sun Jul 10 18:44:55 2022

library IEEE;
use IEEE.std_logic_1164.all;
-- synopsys translate_off
library xp2;
use xp2.components.all;
-- synopsys translate_on

ENTITY byte_cache_16 IS PORT (
   ResetA    : IN  STD_LOGIC;
   ClockA    : IN  STD_LOGIC;
   ClockEnA  : IN  STD_LOGIC;
   WrA       : IN  STD_LOGIC;
   ByteEnA   : IN  STD_LOGIC_VECTOR(1 DOWNTO 0);
   AddressA  : IN  STD_LOGIC_VECTOR(12 DOWNTO 0);
   DataInA   : IN  STD_LOGIC_VECTOR(15 DOWNTO 0);
   QA        : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
-- dma port
   ResetB    : IN  STD_LOGIC;
   ClockB    : IN  STD_LOGIC;
   ClockEnB  : IN  STD_LOGIC;
   WrB       : IN  STD_LOGIC;
   ByteEnB   : IN  STD_LOGIC_VECTOR(1 DOWNTO 0);
   AddressB  : IN  STD_LOGIC_VECTOR(12 DOWNTO 0);
   DataInB   : IN  STD_LOGIC_VECTOR(15 DOWNTO 0);
   QB        : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
); END byte_cache_16;

architecture Structure of byte_cache_16 is

    -- internal signal declarations
    signal scuba_vhi: std_logic;
    signal wren0_inv: std_logic;
    signal wren1_inv: std_logic;
    signal mdout1_0_17: std_logic;
    signal mdout0_0_17: std_logic;
    signal mdout1_0_8: std_logic;
    signal mdout0_0_8: std_logic;
    signal mdout1_1_17: std_logic;
    signal mdout0_1_17: std_logic;
    signal mdout1_1_8: std_logic;
    signal mdout0_1_8: std_logic;
    signal mdout1_2_17: std_logic;
    signal mdout0_2_17: std_logic;
    signal mdout1_2_8: std_logic;
    signal mdout0_2_8: std_logic;
    signal mdout1_3_17: std_logic;
    signal mdout0_3_17: std_logic;
    signal mdout1_3_8: std_logic;
    signal mdout0_3_8: std_logic;
    signal mdout1_4_17: std_logic;
    signal mdout0_4_17: std_logic;
    signal mdout1_4_8: std_logic;
    signal mdout0_4_8: std_logic;
    signal mdout1_5_17: std_logic;
    signal mdout0_5_17: std_logic;
    signal mdout1_5_8: std_logic;
    signal mdout0_5_8: std_logic;
    signal wren0_inv_g: std_logic;
    signal wren1_inv_g: std_logic;
    signal addr110_ff: std_logic;
    signal addr111_ff: std_logic;
    signal addr112_ff: std_logic;
    signal mdout0_5_0: std_logic;
    signal mdout0_4_0: std_logic;
    signal mdout0_3_0: std_logic;
    signal mdout0_2_0: std_logic;
    signal mdout0_1_0: std_logic;
    signal mdout0_0_0: std_logic;
    signal mdout0_5_1: std_logic;
    signal mdout0_4_1: std_logic;
    signal mdout0_3_1: std_logic;
    signal mdout0_2_1: std_logic;
    signal mdout0_1_1: std_logic;
    signal mdout0_0_1: std_logic;
    signal mdout0_5_2: std_logic;
    signal mdout0_4_2: std_logic;
    signal mdout0_3_2: std_logic;
    signal mdout0_2_2: std_logic;
    signal mdout0_1_2: std_logic;
    signal mdout0_0_2: std_logic;
    signal mdout0_5_3: std_logic;
    signal mdout0_4_3: std_logic;
    signal mdout0_3_3: std_logic;
    signal mdout0_2_3: std_logic;
    signal mdout0_1_3: std_logic;
    signal mdout0_0_3: std_logic;
    signal mdout0_5_4: std_logic;
    signal mdout0_4_4: std_logic;
    signal mdout0_3_4: std_logic;
    signal mdout0_2_4: std_logic;
    signal mdout0_1_4: std_logic;
    signal mdout0_0_4: std_logic;
    signal mdout0_5_5: std_logic;
    signal mdout0_4_5: std_logic;
    signal mdout0_3_5: std_logic;
    signal mdout0_2_5: std_logic;
    signal mdout0_1_5: std_logic;
    signal mdout0_0_5: std_logic;
    signal mdout0_5_6: std_logic;
    signal mdout0_4_6: std_logic;
    signal mdout0_3_6: std_logic;
    signal mdout0_2_6: std_logic;
    signal mdout0_1_6: std_logic;
    signal mdout0_0_6: std_logic;
    signal mdout0_5_7: std_logic;
    signal mdout0_4_7: std_logic;
    signal mdout0_3_7: std_logic;
    signal mdout0_2_7: std_logic;
    signal mdout0_1_7: std_logic;
    signal mdout0_0_7: std_logic;
    signal mdout0_5_9: std_logic;
    signal mdout0_4_9: std_logic;
    signal mdout0_3_9: std_logic;
    signal mdout0_2_9: std_logic;
    signal mdout0_1_9: std_logic;
    signal mdout0_0_9: std_logic;
    signal mdout0_5_10: std_logic;
    signal mdout0_4_10: std_logic;
    signal mdout0_3_10: std_logic;
    signal mdout0_2_10: std_logic;
    signal mdout0_1_10: std_logic;
    signal mdout0_0_10: std_logic;
    signal mdout0_5_11: std_logic;
    signal mdout0_4_11: std_logic;
    signal mdout0_3_11: std_logic;
    signal mdout0_2_11: std_logic;
    signal mdout0_1_11: std_logic;
    signal mdout0_0_11: std_logic;
    signal mdout0_5_12: std_logic;
    signal mdout0_4_12: std_logic;
    signal mdout0_3_12: std_logic;
    signal mdout0_2_12: std_logic;
    signal mdout0_1_12: std_logic;
    signal mdout0_0_12: std_logic;
    signal mdout0_5_13: std_logic;
    signal mdout0_4_13: std_logic;
    signal mdout0_3_13: std_logic;
    signal mdout0_2_13: std_logic;
    signal mdout0_1_13: std_logic;
    signal mdout0_0_13: std_logic;
    signal mdout0_5_14: std_logic;
    signal mdout0_4_14: std_logic;
    signal mdout0_3_14: std_logic;
    signal mdout0_2_14: std_logic;
    signal mdout0_1_14: std_logic;
    signal mdout0_0_14: std_logic;
    signal mdout0_5_15: std_logic;
    signal mdout0_4_15: std_logic;
    signal mdout0_3_15: std_logic;
    signal mdout0_2_15: std_logic;
    signal mdout0_1_15: std_logic;
    signal mdout0_0_15: std_logic;
    signal addr012_ff: std_logic;
    signal addr011_ff: std_logic;
    signal addr010_ff: std_logic;
    signal mdout0_5_16: std_logic;
    signal mdout0_4_16: std_logic;
    signal mdout0_3_16: std_logic;
    signal mdout0_2_16: std_logic;
    signal mdout0_1_16: std_logic;
    signal mdout0_0_16: std_logic;
    signal mdout1_5_0: std_logic;
    signal mdout1_4_0: std_logic;
    signal mdout1_3_0: std_logic;
    signal mdout1_2_0: std_logic;
    signal mdout1_1_0: std_logic;
    signal mdout1_0_0: std_logic;
    signal mdout1_5_1: std_logic;
    signal mdout1_4_1: std_logic;
    signal mdout1_3_1: std_logic;
    signal mdout1_2_1: std_logic;
    signal mdout1_1_1: std_logic;
    signal mdout1_0_1: std_logic;
    signal mdout1_5_2: std_logic;
    signal mdout1_4_2: std_logic;
    signal mdout1_3_2: std_logic;
    signal mdout1_2_2: std_logic;
    signal mdout1_1_2: std_logic;
    signal mdout1_0_2: std_logic;
    signal mdout1_5_3: std_logic;
    signal mdout1_4_3: std_logic;
    signal mdout1_3_3: std_logic;
    signal mdout1_2_3: std_logic;
    signal mdout1_1_3: std_logic;
    signal mdout1_0_3: std_logic;
    signal mdout1_5_4: std_logic;
    signal mdout1_4_4: std_logic;
    signal mdout1_3_4: std_logic;
    signal mdout1_2_4: std_logic;
    signal mdout1_1_4: std_logic;
    signal mdout1_0_4: std_logic;
    signal mdout1_5_5: std_logic;
    signal mdout1_4_5: std_logic;
    signal mdout1_3_5: std_logic;
    signal mdout1_2_5: std_logic;
    signal mdout1_1_5: std_logic;
    signal mdout1_0_5: std_logic;
    signal mdout1_5_6: std_logic;
    signal mdout1_4_6: std_logic;
    signal mdout1_3_6: std_logic;
    signal mdout1_2_6: std_logic;
    signal mdout1_1_6: std_logic;
    signal mdout1_0_6: std_logic;
    signal mdout1_5_7: std_logic;
    signal mdout1_4_7: std_logic;
    signal mdout1_3_7: std_logic;
    signal mdout1_2_7: std_logic;
    signal mdout1_1_7: std_logic;
    signal mdout1_0_7: std_logic;
    signal mdout1_5_9: std_logic;
    signal mdout1_4_9: std_logic;
    signal mdout1_3_9: std_logic;
    signal mdout1_2_9: std_logic;
    signal mdout1_1_9: std_logic;
    signal mdout1_0_9: std_logic;
    signal mdout1_5_10: std_logic;
    signal mdout1_4_10: std_logic;
    signal mdout1_3_10: std_logic;
    signal mdout1_2_10: std_logic;
    signal mdout1_1_10: std_logic;
    signal mdout1_0_10: std_logic;
    signal mdout1_5_11: std_logic;
    signal mdout1_4_11: std_logic;
    signal mdout1_3_11: std_logic;
    signal mdout1_2_11: std_logic;
    signal mdout1_1_11: std_logic;
    signal mdout1_0_11: std_logic;
    signal mdout1_5_12: std_logic;
    signal mdout1_4_12: std_logic;
    signal mdout1_3_12: std_logic;
    signal mdout1_2_12: std_logic;
    signal mdout1_1_12: std_logic;
    signal mdout1_0_12: std_logic;
    signal mdout1_5_13: std_logic;
    signal mdout1_4_13: std_logic;
    signal mdout1_3_13: std_logic;
    signal mdout1_2_13: std_logic;
    signal mdout1_1_13: std_logic;
    signal mdout1_0_13: std_logic;
    signal mdout1_5_14: std_logic;
    signal mdout1_4_14: std_logic;
    signal mdout1_3_14: std_logic;
    signal mdout1_2_14: std_logic;
    signal mdout1_1_14: std_logic;
    signal mdout1_0_14: std_logic;
    signal mdout1_5_15: std_logic;
    signal mdout1_4_15: std_logic;
    signal mdout1_3_15: std_logic;
    signal mdout1_2_15: std_logic;
    signal mdout1_1_15: std_logic;
    signal mdout1_0_15: std_logic;
    signal addr112_ff2: std_logic;
    signal addr111_ff2: std_logic;
    signal addr110_ff2: std_logic;
    signal scuba_vlo: std_logic;
    signal mdout1_5_16: std_logic;
    signal mdout1_4_16: std_logic;
    signal mdout1_3_16: std_logic;
    signal mdout1_2_16: std_logic;
    signal mdout1_1_16: std_logic;
    signal mdout1_0_16: std_logic;

    -- local component declarations
    component AND2
        port (A: in  std_logic; B: in  std_logic; Z: out  std_logic);
    end component;
    component FD1P3DX
    -- synopsys translate_off
        generic (GSR : in String);
    -- synopsys translate_on
        port (D: in  std_logic; SP: in  std_logic; CK: in  std_logic;
            CD: in  std_logic; Q: out  std_logic);
    end component;
    component INV
        port (A: in  std_logic; Z: out  std_logic);
    end component;
    component MUX81
        port (D0: in  std_logic; D1: in  std_logic; D2: in  std_logic;
            D3: in  std_logic; D4: in  std_logic; D5: in  std_logic;
            D6: in  std_logic; D7: in  std_logic; SD1: in  std_logic;
            SD2: in  std_logic; SD3: in  std_logic; Z: out  std_logic);
    end component;
    component VHI
        port (Z: out  std_logic);
    end component;
    component VLO
        port (Z: out  std_logic);
    end component;
    component DP16KB
    -- synopsys translate_off
        generic (GSR : in String; WRITEMODE_B : in String;
                CSDECODE_B : in std_logic_vector(2 downto 0);
                CSDECODE_A : in std_logic_vector(2 downto 0);
                WRITEMODE_A : in String; RESETMODE : in String;
                REGMODE_B : in String; REGMODE_A : in String;
                DATA_WIDTH_B : in Integer; DATA_WIDTH_A : in Integer);
    -- synopsys translate_on
        port (DIA0: in  std_logic; DIA1: in  std_logic;
            DIA2: in  std_logic; DIA3: in  std_logic;
            DIA4: in  std_logic; DIA5: in  std_logic;
            DIA6: in  std_logic; DIA7: in  std_logic;
            DIA8: in  std_logic; DIA9: in  std_logic;
            DIA10: in  std_logic; DIA11: in  std_logic;
            DIA12: in  std_logic; DIA13: in  std_logic;
            DIA14: in  std_logic; DIA15: in  std_logic;
            DIA16: in  std_logic; DIA17: in  std_logic;
            ADA0: in  std_logic; ADA1: in  std_logic;
            ADA2: in  std_logic; ADA3: in  std_logic;
            ADA4: in  std_logic; ADA5: in  std_logic;
            ADA6: in  std_logic; ADA7: in  std_logic;
            ADA8: in  std_logic; ADA9: in  std_logic;
            ADA10: in  std_logic; ADA11: in  std_logic;
            ADA12: in  std_logic; ADA13: in  std_logic;
            CEA: in  std_logic; CLKA: in  std_logic; WEA: in  std_logic;
            CSA0: in  std_logic; CSA1: in  std_logic;
            CSA2: in  std_logic; RSTA: in  std_logic;
            DIB0: in  std_logic; DIB1: in  std_logic;
            DIB2: in  std_logic; DIB3: in  std_logic;
            DIB4: in  std_logic; DIB5: in  std_logic;
            DIB6: in  std_logic; DIB7: in  std_logic;
            DIB8: in  std_logic; DIB9: in  std_logic;
            DIB10: in  std_logic; DIB11: in  std_logic;
            DIB12: in  std_logic; DIB13: in  std_logic;
            DIB14: in  std_logic; DIB15: in  std_logic;
            DIB16: in  std_logic; DIB17: in  std_logic;
            ADB0: in  std_logic; ADB1: in  std_logic;
            ADB2: in  std_logic; ADB3: in  std_logic;
            ADB4: in  std_logic; ADB5: in  std_logic;
            ADB6: in  std_logic; ADB7: in  std_logic;
            ADB8: in  std_logic; ADB9: in  std_logic;
            ADB10: in  std_logic; ADB11: in  std_logic;
            ADB12: in  std_logic; ADB13: in  std_logic;
            CEB: in  std_logic; CLKB: in  std_logic; WEB: in  std_logic;
            CSB0: in  std_logic; CSB1: in  std_logic;
            CSB2: in  std_logic; RSTB: in  std_logic;
            DOA0: out  std_logic; DOA1: out  std_logic;
            DOA2: out  std_logic; DOA3: out  std_logic;
            DOA4: out  std_logic; DOA5: out  std_logic;
            DOA6: out  std_logic; DOA7: out  std_logic;
            DOA8: out  std_logic; DOA9: out  std_logic;
            DOA10: out  std_logic; DOA11: out  std_logic;
            DOA12: out  std_logic; DOA13: out  std_logic;
            DOA14: out  std_logic; DOA15: out  std_logic;
            DOA16: out  std_logic; DOA17: out  std_logic;
            DOB0: out  std_logic; DOB1: out  std_logic;
            DOB2: out  std_logic; DOB3: out  std_logic;
            DOB4: out  std_logic; DOB5: out  std_logic;
            DOB6: out  std_logic; DOB7: out  std_logic;
            DOB8: out  std_logic; DOB9: out  std_logic;
            DOB10: out  std_logic; DOB11: out  std_logic;
            DOB12: out  std_logic; DOB13: out  std_logic;
            DOB14: out  std_logic; DOB15: out  std_logic;
            DOB16: out  std_logic; DOB17: out  std_logic);
    end component;
    attribute MEM_LPC_FILE : string;
    attribute MEM_INIT_FILE : string;
    attribute CSDECODE_B : string;
    attribute CSDECODE_A : string;
    attribute WRITEMODE_B : string;
    attribute WRITEMODE_A : string;
    attribute RESETMODE : string;
    attribute REGMODE_B : string;
    attribute REGMODE_A : string;
    attribute DATA_WIDTH_B : string;
    attribute DATA_WIDTH_A : string;
    attribute GSR : string;
    attribute MEM_LPC_FILE of byte_cache_16_0_0_5 : label is "byte_cache_16.lpc";
    attribute MEM_INIT_FILE of byte_cache_16_0_0_5 : label is "";
    attribute CSDECODE_B of byte_cache_16_0_0_5 : label is "0b000";
    attribute CSDECODE_A of byte_cache_16_0_0_5 : label is "0b000";
    attribute WRITEMODE_B of byte_cache_16_0_0_5 : label is "NORMAL";
    attribute WRITEMODE_A of byte_cache_16_0_0_5 : label is "NORMAL";
    attribute GSR of byte_cache_16_0_0_5 : label is "DISABLED";
    attribute RESETMODE of byte_cache_16_0_0_5 : label is "SYNC";
    attribute REGMODE_B of byte_cache_16_0_0_5 : label is "OUTREG";
    attribute REGMODE_A of byte_cache_16_0_0_5 : label is "NOREG";
    attribute DATA_WIDTH_B of byte_cache_16_0_0_5 : label is "18";
    attribute DATA_WIDTH_A of byte_cache_16_0_0_5 : label is "18";
    attribute MEM_LPC_FILE of byte_cache_16_1_0_4 : label is "byte_cache_16.lpc";
    attribute MEM_INIT_FILE of byte_cache_16_1_0_4 : label is "";
    attribute CSDECODE_B of byte_cache_16_1_0_4 : label is "0b001";
    attribute CSDECODE_A of byte_cache_16_1_0_4 : label is "0b001";
    attribute WRITEMODE_B of byte_cache_16_1_0_4 : label is "NORMAL";
    attribute WRITEMODE_A of byte_cache_16_1_0_4 : label is "NORMAL";
    attribute GSR of byte_cache_16_1_0_4 : label is "DISABLED";
    attribute RESETMODE of byte_cache_16_1_0_4 : label is "SYNC";
    attribute REGMODE_B of byte_cache_16_1_0_4 : label is "OUTREG";
    attribute REGMODE_A of byte_cache_16_1_0_4 : label is "NOREG";
    attribute DATA_WIDTH_B of byte_cache_16_1_0_4 : label is "18";
    attribute DATA_WIDTH_A of byte_cache_16_1_0_4 : label is "18";
    attribute MEM_LPC_FILE of byte_cache_16_2_0_3 : label is "byte_cache_16.lpc";
    attribute MEM_INIT_FILE of byte_cache_16_2_0_3 : label is "";
    attribute CSDECODE_B of byte_cache_16_2_0_3 : label is "0b010";
    attribute CSDECODE_A of byte_cache_16_2_0_3 : label is "0b010";
    attribute WRITEMODE_B of byte_cache_16_2_0_3 : label is "NORMAL";
    attribute WRITEMODE_A of byte_cache_16_2_0_3 : label is "NORMAL";
    attribute GSR of byte_cache_16_2_0_3 : label is "DISABLED";
    attribute RESETMODE of byte_cache_16_2_0_3 : label is "SYNC";
    attribute REGMODE_B of byte_cache_16_2_0_3 : label is "OUTREG";
    attribute REGMODE_A of byte_cache_16_2_0_3 : label is "NOREG";
    attribute DATA_WIDTH_B of byte_cache_16_2_0_3 : label is "18";
    attribute DATA_WIDTH_A of byte_cache_16_2_0_3 : label is "18";
    attribute MEM_LPC_FILE of byte_cache_16_3_0_2 : label is "byte_cache_16.lpc";
    attribute MEM_INIT_FILE of byte_cache_16_3_0_2 : label is "";
    attribute CSDECODE_B of byte_cache_16_3_0_2 : label is "0b011";
    attribute CSDECODE_A of byte_cache_16_3_0_2 : label is "0b011";
    attribute WRITEMODE_B of byte_cache_16_3_0_2 : label is "NORMAL";
    attribute WRITEMODE_A of byte_cache_16_3_0_2 : label is "NORMAL";
    attribute GSR of byte_cache_16_3_0_2 : label is "DISABLED";
    attribute RESETMODE of byte_cache_16_3_0_2 : label is "SYNC";
    attribute REGMODE_B of byte_cache_16_3_0_2 : label is "OUTREG";
    attribute REGMODE_A of byte_cache_16_3_0_2 : label is "NOREG";
    attribute DATA_WIDTH_B of byte_cache_16_3_0_2 : label is "18";
    attribute DATA_WIDTH_A of byte_cache_16_3_0_2 : label is "18";
    attribute MEM_LPC_FILE of byte_cache_16_4_0_1 : label is "byte_cache_16.lpc";
    attribute MEM_INIT_FILE of byte_cache_16_4_0_1 : label is "";
    attribute CSDECODE_B of byte_cache_16_4_0_1 : label is "0b100";
    attribute CSDECODE_A of byte_cache_16_4_0_1 : label is "0b100";
    attribute WRITEMODE_B of byte_cache_16_4_0_1 : label is "NORMAL";
    attribute WRITEMODE_A of byte_cache_16_4_0_1 : label is "NORMAL";
    attribute GSR of byte_cache_16_4_0_1 : label is "DISABLED";
    attribute RESETMODE of byte_cache_16_4_0_1 : label is "SYNC";
    attribute REGMODE_B of byte_cache_16_4_0_1 : label is "OUTREG";
    attribute REGMODE_A of byte_cache_16_4_0_1 : label is "NOREG";
    attribute DATA_WIDTH_B of byte_cache_16_4_0_1 : label is "18";
    attribute DATA_WIDTH_A of byte_cache_16_4_0_1 : label is "18";
    attribute MEM_LPC_FILE of byte_cache_16_5_0_0 : label is "byte_cache_16.lpc";
    attribute MEM_INIT_FILE of byte_cache_16_5_0_0 : label is "";
    attribute CSDECODE_B of byte_cache_16_5_0_0 : label is "0b101";
    attribute CSDECODE_A of byte_cache_16_5_0_0 : label is "0b101";
    attribute WRITEMODE_B of byte_cache_16_5_0_0 : label is "NORMAL";
    attribute WRITEMODE_A of byte_cache_16_5_0_0 : label is "NORMAL";
    attribute GSR of byte_cache_16_5_0_0 : label is "DISABLED";
    attribute RESETMODE of byte_cache_16_5_0_0 : label is "SYNC";
    attribute REGMODE_B of byte_cache_16_5_0_0 : label is "OUTREG";
    attribute REGMODE_A of byte_cache_16_5_0_0 : label is "NOREG";
    attribute DATA_WIDTH_B of byte_cache_16_5_0_0 : label is "18";
    attribute DATA_WIDTH_A of byte_cache_16_5_0_0 : label is "18";
    attribute GSR of FF_8 : label is "ENABLED";
    attribute GSR of FF_7 : label is "ENABLED";
    attribute GSR of FF_6 : label is "ENABLED";
    attribute GSR of FF_5 : label is "ENABLED";
    attribute GSR of FF_4 : label is "ENABLED";
    attribute GSR of FF_3 : label is "ENABLED";
    attribute GSR of FF_2 : label is "ENABLED";
    attribute GSR of FF_1 : label is "ENABLED";
    attribute GSR of FF_0 : label is "ENABLED";
    attribute NGD_DRC_MASK : integer;
    attribute NGD_DRC_MASK of Structure : architecture is 1;

begin
    -- component instantiation statements
    scuba_vhi_inst: VHI
        port map (Z=>scuba_vhi);

    INV_1: INV
        port map (A=>WrA, Z=>wren0_inv);

    AND2_t1: AND2
        port map (A=>wren0_inv, B=>ClockEnA, Z=>wren0_inv_g);

    INV_0: INV
        port map (A=>WrB, Z=>wren1_inv);

    AND2_t0: AND2
        port map (A=>wren1_inv, B=>ClockEnB, Z=>wren1_inv_g);

    byte_cache_16_0_0_5: DP16KB
        -- synopsys translate_off
        generic map (CSDECODE_B=> "000", CSDECODE_A=> "000", WRITEMODE_B=> "NORMAL",
        WRITEMODE_A=> "NORMAL", GSR=> "DISABLED", RESETMODE=> "SYNC",
        REGMODE_B=> "OUTREG", REGMODE_A=> "NOREG", DATA_WIDTH_B=>  18,
        DATA_WIDTH_A=>  18)
        -- synopsys translate_on
        port map (DIA0=>DataInA(0), DIA1=>DataInA(1), DIA2=>DataInA(2),
            DIA3=>DataInA(3), DIA4=>DataInA(4), DIA5=>DataInA(5),
            DIA6=>DataInA(6), DIA7=>DataInA(7), DIA8=>scuba_vlo,
            DIA9=>DataInA(8), DIA10=>DataInA(9), DIA11=>DataInA(10),
            DIA12=>DataInA(11), DIA13=>DataInA(12), DIA14=>DataInA(13),
            DIA15=>DataInA(14), DIA16=>DataInA(15), DIA17=>scuba_vlo,
            ADA0=>ByteEnA(0), ADA1=>ByteEnA(1), ADA2=>scuba_vlo,
            ADA3=>scuba_vlo, ADA4=>AddressA(0), ADA5=>AddressA(1),
            ADA6=>AddressA(2), ADA7=>AddressA(3), ADA8=>AddressA(4),
            ADA9=>AddressA(5), ADA10=>AddressA(6), ADA11=>AddressA(7),
            ADA12=>AddressA(8), ADA13=>AddressA(9), CEA=>ClockEnA,
            CLKA=>ClockA, WEA=>WrA, CSA0=>AddressA(10),
            CSA1=>AddressA(11), CSA2=>AddressA(12), RSTA=>ResetA,
            DIB0=>DataInB(0), DIB1=>DataInB(1), DIB2=>DataInB(2),
            DIB3=>DataInB(3), DIB4=>DataInB(4), DIB5=>DataInB(5),
            DIB6=>DataInB(6), DIB7=>DataInB(7), DIB8=>scuba_vlo,
            DIB9=>DataInB(8), DIB10=>DataInB(9), DIB11=>DataInB(10),
            DIB12=>DataInB(11), DIB13=>DataInB(12), DIB14=>DataInB(13),
            DIB15=>DataInB(14), DIB16=>DataInB(15), DIB17=>scuba_vlo,
            ADB0=>ByteEnB(0), ADB1=>ByteEnB(1), ADB2=>scuba_vlo,
            ADB3=>scuba_vlo, ADB4=>AddressB(0), ADB5=>AddressB(1),
            ADB6=>AddressB(2), ADB7=>AddressB(3), ADB8=>AddressB(4),
            ADB9=>AddressB(5), ADB10=>AddressB(6), ADB11=>AddressB(7),
            ADB12=>AddressB(8), ADB13=>AddressB(9), CEB=>ClockEnB,
            CLKB=>ClockB, WEB=>WrB, CSB0=>AddressB(10),
            CSB1=>AddressB(11), CSB2=>AddressB(12), RSTB=>ResetB,
            DOA0=>mdout0_0_0, DOA1=>mdout0_0_1, DOA2=>mdout0_0_2,
            DOA3=>mdout0_0_3, DOA4=>mdout0_0_4, DOA5=>mdout0_0_5,
            DOA6=>mdout0_0_6, DOA7=>mdout0_0_7, DOA8=>mdout0_0_8,
            DOA9=>mdout0_0_9, DOA10=>mdout0_0_10, DOA11=>mdout0_0_11,
            DOA12=>mdout0_0_12, DOA13=>mdout0_0_13, DOA14=>mdout0_0_14,
            DOA15=>mdout0_0_15, DOA16=>mdout0_0_16, DOA17=>mdout0_0_17,
            DOB0=>mdout1_0_0, DOB1=>mdout1_0_1, DOB2=>mdout1_0_2,
            DOB3=>mdout1_0_3, DOB4=>mdout1_0_4, DOB5=>mdout1_0_5,
            DOB6=>mdout1_0_6, DOB7=>mdout1_0_7, DOB8=>mdout1_0_8,
            DOB9=>mdout1_0_9, DOB10=>mdout1_0_10, DOB11=>mdout1_0_11,
            DOB12=>mdout1_0_12, DOB13=>mdout1_0_13, DOB14=>mdout1_0_14,
            DOB15=>mdout1_0_15, DOB16=>mdout1_0_16, DOB17=>mdout1_0_17);

    byte_cache_16_1_0_4: DP16KB
        -- synopsys translate_off
        generic map (CSDECODE_B=> "001", CSDECODE_A=> "001", WRITEMODE_B=> "NORMAL",
        WRITEMODE_A=> "NORMAL", GSR=> "DISABLED", RESETMODE=> "SYNC",
        REGMODE_B=> "OUTREG", REGMODE_A=> "NOREG", DATA_WIDTH_B=>  18,
        DATA_WIDTH_A=>  18)
        -- synopsys translate_on
        port map (DIA0=>DataInA(0), DIA1=>DataInA(1), DIA2=>DataInA(2),
            DIA3=>DataInA(3), DIA4=>DataInA(4), DIA5=>DataInA(5),
            DIA6=>DataInA(6), DIA7=>DataInA(7), DIA8=>scuba_vlo,
            DIA9=>DataInA(8), DIA10=>DataInA(9), DIA11=>DataInA(10),
            DIA12=>DataInA(11), DIA13=>DataInA(12), DIA14=>DataInA(13),
            DIA15=>DataInA(14), DIA16=>DataInA(15), DIA17=>scuba_vlo,
            ADA0=>ByteEnA(0), ADA1=>ByteEnA(1), ADA2=>scuba_vlo,
            ADA3=>scuba_vlo, ADA4=>AddressA(0), ADA5=>AddressA(1),
            ADA6=>AddressA(2), ADA7=>AddressA(3), ADA8=>AddressA(4),
            ADA9=>AddressA(5), ADA10=>AddressA(6), ADA11=>AddressA(7),
            ADA12=>AddressA(8), ADA13=>AddressA(9), CEA=>ClockEnA,
            CLKA=>ClockA, WEA=>WrA, CSA0=>AddressA(10),
            CSA1=>AddressA(11), CSA2=>AddressA(12), RSTA=>ResetA,
            DIB0=>DataInB(0), DIB1=>DataInB(1), DIB2=>DataInB(2),
            DIB3=>DataInB(3), DIB4=>DataInB(4), DIB5=>DataInB(5),
            DIB6=>DataInB(6), DIB7=>DataInB(7), DIB8=>scuba_vlo,
            DIB9=>DataInB(8), DIB10=>DataInB(9), DIB11=>DataInB(10),
            DIB12=>DataInB(11), DIB13=>DataInB(12), DIB14=>DataInB(13),
            DIB15=>DataInB(14), DIB16=>DataInB(15), DIB17=>scuba_vlo,
            ADB0=>ByteEnB(0), ADB1=>ByteEnB(1), ADB2=>scuba_vlo,
            ADB3=>scuba_vlo, ADB4=>AddressB(0), ADB5=>AddressB(1),
            ADB6=>AddressB(2), ADB7=>AddressB(3), ADB8=>AddressB(4),
            ADB9=>AddressB(5), ADB10=>AddressB(6), ADB11=>AddressB(7),
            ADB12=>AddressB(8), ADB13=>AddressB(9), CEB=>ClockEnB,
            CLKB=>ClockB, WEB=>WrB, CSB0=>AddressB(10),
            CSB1=>AddressB(11), CSB2=>AddressB(12), RSTB=>ResetB,
            DOA0=>mdout0_1_0, DOA1=>mdout0_1_1, DOA2=>mdout0_1_2,
            DOA3=>mdout0_1_3, DOA4=>mdout0_1_4, DOA5=>mdout0_1_5,
            DOA6=>mdout0_1_6, DOA7=>mdout0_1_7, DOA8=>mdout0_1_8,
            DOA9=>mdout0_1_9, DOA10=>mdout0_1_10, DOA11=>mdout0_1_11,
            DOA12=>mdout0_1_12, DOA13=>mdout0_1_13, DOA14=>mdout0_1_14,
            DOA15=>mdout0_1_15, DOA16=>mdout0_1_16, DOA17=>mdout0_1_17,
            DOB0=>mdout1_1_0, DOB1=>mdout1_1_1, DOB2=>mdout1_1_2,
            DOB3=>mdout1_1_3, DOB4=>mdout1_1_4, DOB5=>mdout1_1_5,
            DOB6=>mdout1_1_6, DOB7=>mdout1_1_7, DOB8=>mdout1_1_8,
            DOB9=>mdout1_1_9, DOB10=>mdout1_1_10, DOB11=>mdout1_1_11,
            DOB12=>mdout1_1_12, DOB13=>mdout1_1_13, DOB14=>mdout1_1_14,
            DOB15=>mdout1_1_15, DOB16=>mdout1_1_16, DOB17=>mdout1_1_17);

    byte_cache_16_2_0_3: DP16KB
        -- synopsys translate_off
        generic map (CSDECODE_B=> "010", CSDECODE_A=> "010", WRITEMODE_B=> "NORMAL",
        WRITEMODE_A=> "NORMAL", GSR=> "DISABLED", RESETMODE=> "SYNC",
        REGMODE_B=> "OUTREG", REGMODE_A=> "NOREG", DATA_WIDTH_B=>  18,
        DATA_WIDTH_A=>  18)
        -- synopsys translate_on
        port map (DIA0=>DataInA(0), DIA1=>DataInA(1), DIA2=>DataInA(2),
            DIA3=>DataInA(3), DIA4=>DataInA(4), DIA5=>DataInA(5),
            DIA6=>DataInA(6), DIA7=>DataInA(7), DIA8=>scuba_vlo,
            DIA9=>DataInA(8), DIA10=>DataInA(9), DIA11=>DataInA(10),
            DIA12=>DataInA(11), DIA13=>DataInA(12), DIA14=>DataInA(13),
            DIA15=>DataInA(14), DIA16=>DataInA(15), DIA17=>scuba_vlo,
            ADA0=>ByteEnA(0), ADA1=>ByteEnA(1), ADA2=>scuba_vlo,
            ADA3=>scuba_vlo, ADA4=>AddressA(0), ADA5=>AddressA(1),
            ADA6=>AddressA(2), ADA7=>AddressA(3), ADA8=>AddressA(4),
            ADA9=>AddressA(5), ADA10=>AddressA(6), ADA11=>AddressA(7),
            ADA12=>AddressA(8), ADA13=>AddressA(9), CEA=>ClockEnA,
            CLKA=>ClockA, WEA=>WrA, CSA0=>AddressA(10),
            CSA1=>AddressA(11), CSA2=>AddressA(12), RSTA=>ResetA,
            DIB0=>DataInB(0), DIB1=>DataInB(1), DIB2=>DataInB(2),
            DIB3=>DataInB(3), DIB4=>DataInB(4), DIB5=>DataInB(5),
            DIB6=>DataInB(6), DIB7=>DataInB(7), DIB8=>scuba_vlo,
            DIB9=>DataInB(8), DIB10=>DataInB(9), DIB11=>DataInB(10),
            DIB12=>DataInB(11), DIB13=>DataInB(12), DIB14=>DataInB(13),
            DIB15=>DataInB(14), DIB16=>DataInB(15), DIB17=>scuba_vlo,
            ADB0=>ByteEnB(0), ADB1=>ByteEnB(1), ADB2=>scuba_vlo,
            ADB3=>scuba_vlo, ADB4=>AddressB(0), ADB5=>AddressB(1),
            ADB6=>AddressB(2), ADB7=>AddressB(3), ADB8=>AddressB(4),
            ADB9=>AddressB(5), ADB10=>AddressB(6), ADB11=>AddressB(7),
            ADB12=>AddressB(8), ADB13=>AddressB(9), CEB=>ClockEnB,
            CLKB=>ClockB, WEB=>WrB, CSB0=>AddressB(10),
            CSB1=>AddressB(11), CSB2=>AddressB(12), RSTB=>ResetB,
            DOA0=>mdout0_2_0, DOA1=>mdout0_2_1, DOA2=>mdout0_2_2,
            DOA3=>mdout0_2_3, DOA4=>mdout0_2_4, DOA5=>mdout0_2_5,
            DOA6=>mdout0_2_6, DOA7=>mdout0_2_7, DOA8=>mdout0_2_8,
            DOA9=>mdout0_2_9, DOA10=>mdout0_2_10, DOA11=>mdout0_2_11,
            DOA12=>mdout0_2_12, DOA13=>mdout0_2_13, DOA14=>mdout0_2_14,
            DOA15=>mdout0_2_15, DOA16=>mdout0_2_16, DOA17=>mdout0_2_17,
            DOB0=>mdout1_2_0, DOB1=>mdout1_2_1, DOB2=>mdout1_2_2,
            DOB3=>mdout1_2_3, DOB4=>mdout1_2_4, DOB5=>mdout1_2_5,
            DOB6=>mdout1_2_6, DOB7=>mdout1_2_7, DOB8=>mdout1_2_8,
            DOB9=>mdout1_2_9, DOB10=>mdout1_2_10, DOB11=>mdout1_2_11,
            DOB12=>mdout1_2_12, DOB13=>mdout1_2_13, DOB14=>mdout1_2_14,
            DOB15=>mdout1_2_15, DOB16=>mdout1_2_16, DOB17=>mdout1_2_17);

    byte_cache_16_3_0_2: DP16KB
        -- synopsys translate_off
        generic map (CSDECODE_B=> "011", CSDECODE_A=> "011", WRITEMODE_B=> "NORMAL",
        WRITEMODE_A=> "NORMAL", GSR=> "DISABLED", RESETMODE=> "SYNC",
        REGMODE_B=> "OUTREG", REGMODE_A=> "NOREG", DATA_WIDTH_B=>  18,
        DATA_WIDTH_A=>  18)
        -- synopsys translate_on
        port map (DIA0=>DataInA(0), DIA1=>DataInA(1), DIA2=>DataInA(2),
            DIA3=>DataInA(3), DIA4=>DataInA(4), DIA5=>DataInA(5),
            DIA6=>DataInA(6), DIA7=>DataInA(7), DIA8=>scuba_vlo,
            DIA9=>DataInA(8), DIA10=>DataInA(9), DIA11=>DataInA(10),
            DIA12=>DataInA(11), DIA13=>DataInA(12), DIA14=>DataInA(13),
            DIA15=>DataInA(14), DIA16=>DataInA(15), DIA17=>scuba_vlo,
            ADA0=>ByteEnA(0), ADA1=>ByteEnA(1), ADA2=>scuba_vlo,
            ADA3=>scuba_vlo, ADA4=>AddressA(0), ADA5=>AddressA(1),
            ADA6=>AddressA(2), ADA7=>AddressA(3), ADA8=>AddressA(4),
            ADA9=>AddressA(5), ADA10=>AddressA(6), ADA11=>AddressA(7),
            ADA12=>AddressA(8), ADA13=>AddressA(9), CEA=>ClockEnA,
            CLKA=>ClockA, WEA=>WrA, CSA0=>AddressA(10),
            CSA1=>AddressA(11), CSA2=>AddressA(12), RSTA=>ResetA,
            DIB0=>DataInB(0), DIB1=>DataInB(1), DIB2=>DataInB(2),
            DIB3=>DataInB(3), DIB4=>DataInB(4), DIB5=>DataInB(5),
            DIB6=>DataInB(6), DIB7=>DataInB(7), DIB8=>scuba_vlo,
            DIB9=>DataInB(8), DIB10=>DataInB(9), DIB11=>DataInB(10),
            DIB12=>DataInB(11), DIB13=>DataInB(12), DIB14=>DataInB(13),
            DIB15=>DataInB(14), DIB16=>DataInB(15), DIB17=>scuba_vlo,
            ADB0=>ByteEnB(0), ADB1=>ByteEnB(1), ADB2=>scuba_vlo,
            ADB3=>scuba_vlo, ADB4=>AddressB(0), ADB5=>AddressB(1),
            ADB6=>AddressB(2), ADB7=>AddressB(3), ADB8=>AddressB(4),
            ADB9=>AddressB(5), ADB10=>AddressB(6), ADB11=>AddressB(7),
            ADB12=>AddressB(8), ADB13=>AddressB(9), CEB=>ClockEnB,
            CLKB=>ClockB, WEB=>WrB, CSB0=>AddressB(10),
            CSB1=>AddressB(11), CSB2=>AddressB(12), RSTB=>ResetB,
            DOA0=>mdout0_3_0, DOA1=>mdout0_3_1, DOA2=>mdout0_3_2,
            DOA3=>mdout0_3_3, DOA4=>mdout0_3_4, DOA5=>mdout0_3_5,
            DOA6=>mdout0_3_6, DOA7=>mdout0_3_7, DOA8=>mdout0_3_8,
            DOA9=>mdout0_3_9, DOA10=>mdout0_3_10, DOA11=>mdout0_3_11,
            DOA12=>mdout0_3_12, DOA13=>mdout0_3_13, DOA14=>mdout0_3_14,
            DOA15=>mdout0_3_15, DOA16=>mdout0_3_16, DOA17=>mdout0_3_17,
            DOB0=>mdout1_3_0, DOB1=>mdout1_3_1, DOB2=>mdout1_3_2,
            DOB3=>mdout1_3_3, DOB4=>mdout1_3_4, DOB5=>mdout1_3_5,
            DOB6=>mdout1_3_6, DOB7=>mdout1_3_7, DOB8=>mdout1_3_8,
            DOB9=>mdout1_3_9, DOB10=>mdout1_3_10, DOB11=>mdout1_3_11,
            DOB12=>mdout1_3_12, DOB13=>mdout1_3_13, DOB14=>mdout1_3_14,
            DOB15=>mdout1_3_15, DOB16=>mdout1_3_16, DOB17=>mdout1_3_17);

    byte_cache_16_4_0_1: DP16KB
        -- synopsys translate_off
        generic map (CSDECODE_B=> "100", CSDECODE_A=> "100", WRITEMODE_B=> "NORMAL",
        WRITEMODE_A=> "NORMAL", GSR=> "DISABLED", RESETMODE=> "SYNC",
        REGMODE_B=> "OUTREG", REGMODE_A=> "NOREG", DATA_WIDTH_B=>  18,
        DATA_WIDTH_A=>  18)
        -- synopsys translate_on
        port map (DIA0=>DataInA(0), DIA1=>DataInA(1), DIA2=>DataInA(2),
            DIA3=>DataInA(3), DIA4=>DataInA(4), DIA5=>DataInA(5),
            DIA6=>DataInA(6), DIA7=>DataInA(7), DIA8=>scuba_vlo,
            DIA9=>DataInA(8), DIA10=>DataInA(9), DIA11=>DataInA(10),
            DIA12=>DataInA(11), DIA13=>DataInA(12), DIA14=>DataInA(13),
            DIA15=>DataInA(14), DIA16=>DataInA(15), DIA17=>scuba_vlo,
            ADA0=>ByteEnA(0), ADA1=>ByteEnA(1), ADA2=>scuba_vlo,
            ADA3=>scuba_vlo, ADA4=>AddressA(0), ADA5=>AddressA(1),
            ADA6=>AddressA(2), ADA7=>AddressA(3), ADA8=>AddressA(4),
            ADA9=>AddressA(5), ADA10=>AddressA(6), ADA11=>AddressA(7),
            ADA12=>AddressA(8), ADA13=>AddressA(9), CEA=>ClockEnA,
            CLKA=>ClockA, WEA=>WrA, CSA0=>AddressA(10),
            CSA1=>AddressA(11), CSA2=>AddressA(12), RSTA=>ResetA,
            DIB0=>DataInB(0), DIB1=>DataInB(1), DIB2=>DataInB(2),
            DIB3=>DataInB(3), DIB4=>DataInB(4), DIB5=>DataInB(5),
            DIB6=>DataInB(6), DIB7=>DataInB(7), DIB8=>scuba_vlo,
            DIB9=>DataInB(8), DIB10=>DataInB(9), DIB11=>DataInB(10),
            DIB12=>DataInB(11), DIB13=>DataInB(12), DIB14=>DataInB(13),
            DIB15=>DataInB(14), DIB16=>DataInB(15), DIB17=>scuba_vlo,
            ADB0=>ByteEnB(0), ADB1=>ByteEnB(1), ADB2=>scuba_vlo,
            ADB3=>scuba_vlo, ADB4=>AddressB(0), ADB5=>AddressB(1),
            ADB6=>AddressB(2), ADB7=>AddressB(3), ADB8=>AddressB(4),
            ADB9=>AddressB(5), ADB10=>AddressB(6), ADB11=>AddressB(7),
            ADB12=>AddressB(8), ADB13=>AddressB(9), CEB=>ClockEnB,
            CLKB=>ClockB, WEB=>WrB, CSB0=>AddressB(10),
            CSB1=>AddressB(11), CSB2=>AddressB(12), RSTB=>ResetB,
            DOA0=>mdout0_4_0, DOA1=>mdout0_4_1, DOA2=>mdout0_4_2,
            DOA3=>mdout0_4_3, DOA4=>mdout0_4_4, DOA5=>mdout0_4_5,
            DOA6=>mdout0_4_6, DOA7=>mdout0_4_7, DOA8=>mdout0_4_8,
            DOA9=>mdout0_4_9, DOA10=>mdout0_4_10, DOA11=>mdout0_4_11,
            DOA12=>mdout0_4_12, DOA13=>mdout0_4_13, DOA14=>mdout0_4_14,
            DOA15=>mdout0_4_15, DOA16=>mdout0_4_16, DOA17=>mdout0_4_17,
            DOB0=>mdout1_4_0, DOB1=>mdout1_4_1, DOB2=>mdout1_4_2,
            DOB3=>mdout1_4_3, DOB4=>mdout1_4_4, DOB5=>mdout1_4_5,
            DOB6=>mdout1_4_6, DOB7=>mdout1_4_7, DOB8=>mdout1_4_8,
            DOB9=>mdout1_4_9, DOB10=>mdout1_4_10, DOB11=>mdout1_4_11,
            DOB12=>mdout1_4_12, DOB13=>mdout1_4_13, DOB14=>mdout1_4_14,
            DOB15=>mdout1_4_15, DOB16=>mdout1_4_16, DOB17=>mdout1_4_17);

    byte_cache_16_5_0_0: DP16KB
        -- synopsys translate_off
        generic map (CSDECODE_B=> "101", CSDECODE_A=> "101", WRITEMODE_B=> "NORMAL",
        WRITEMODE_A=> "NORMAL", GSR=> "DISABLED", RESETMODE=> "SYNC",
        REGMODE_B=> "OUTREG", REGMODE_A=> "NOREG", DATA_WIDTH_B=>  18,
        DATA_WIDTH_A=>  18)
        -- synopsys translate_on
        port map (DIA0=>DataInA(0), DIA1=>DataInA(1), DIA2=>DataInA(2),
            DIA3=>DataInA(3), DIA4=>DataInA(4), DIA5=>DataInA(5),
            DIA6=>DataInA(6), DIA7=>DataInA(7), DIA8=>scuba_vlo,
            DIA9=>DataInA(8), DIA10=>DataInA(9), DIA11=>DataInA(10),
            DIA12=>DataInA(11), DIA13=>DataInA(12), DIA14=>DataInA(13),
            DIA15=>DataInA(14), DIA16=>DataInA(15), DIA17=>scuba_vlo,
            ADA0=>ByteEnA(0), ADA1=>ByteEnA(1), ADA2=>scuba_vlo,
            ADA3=>scuba_vlo, ADA4=>AddressA(0), ADA5=>AddressA(1),
            ADA6=>AddressA(2), ADA7=>AddressA(3), ADA8=>AddressA(4),
            ADA9=>AddressA(5), ADA10=>AddressA(6), ADA11=>AddressA(7),
            ADA12=>AddressA(8), ADA13=>AddressA(9), CEA=>ClockEnA,
            CLKA=>ClockA, WEA=>WrA, CSA0=>AddressA(10),
            CSA1=>AddressA(11), CSA2=>AddressA(12), RSTA=>ResetA,
            DIB0=>DataInB(0), DIB1=>DataInB(1), DIB2=>DataInB(2),
            DIB3=>DataInB(3), DIB4=>DataInB(4), DIB5=>DataInB(5),
            DIB6=>DataInB(6), DIB7=>DataInB(7), DIB8=>scuba_vlo,
            DIB9=>DataInB(8), DIB10=>DataInB(9), DIB11=>DataInB(10),
            DIB12=>DataInB(11), DIB13=>DataInB(12), DIB14=>DataInB(13),
            DIB15=>DataInB(14), DIB16=>DataInB(15), DIB17=>scuba_vlo,
            ADB0=>ByteEnB(0), ADB1=>ByteEnB(1), ADB2=>scuba_vlo,
            ADB3=>scuba_vlo, ADB4=>AddressB(0), ADB5=>AddressB(1),
            ADB6=>AddressB(2), ADB7=>AddressB(3), ADB8=>AddressB(4),
            ADB9=>AddressB(5), ADB10=>AddressB(6), ADB11=>AddressB(7),
            ADB12=>AddressB(8), ADB13=>AddressB(9), CEB=>ClockEnB,
            CLKB=>ClockB, WEB=>WrB, CSB0=>AddressB(10),
            CSB1=>AddressB(11), CSB2=>AddressB(12), RSTB=>ResetB,
            DOA0=>mdout0_5_0, DOA1=>mdout0_5_1, DOA2=>mdout0_5_2,
            DOA3=>mdout0_5_3, DOA4=>mdout0_5_4, DOA5=>mdout0_5_5,
            DOA6=>mdout0_5_6, DOA7=>mdout0_5_7, DOA8=>mdout0_5_8,
            DOA9=>mdout0_5_9, DOA10=>mdout0_5_10, DOA11=>mdout0_5_11,
            DOA12=>mdout0_5_12, DOA13=>mdout0_5_13, DOA14=>mdout0_5_14,
            DOA15=>mdout0_5_15, DOA16=>mdout0_5_16, DOA17=>mdout0_5_17,
            DOB0=>mdout1_5_0, DOB1=>mdout1_5_1, DOB2=>mdout1_5_2,
            DOB3=>mdout1_5_3, DOB4=>mdout1_5_4, DOB5=>mdout1_5_5,
            DOB6=>mdout1_5_6, DOB7=>mdout1_5_7, DOB8=>mdout1_5_8,
            DOB9=>mdout1_5_9, DOB10=>mdout1_5_10, DOB11=>mdout1_5_11,
            DOB12=>mdout1_5_12, DOB13=>mdout1_5_13, DOB14=>mdout1_5_14,
            DOB15=>mdout1_5_15, DOB16=>mdout1_5_16, DOB17=>mdout1_5_17);

    FF_8: FD1P3DX
        -- synopsys translate_off
        generic map (GSR=> "ENABLED")
        -- synopsys translate_on
        port map (D=>AddressA(10), SP=>wren0_inv_g, CK=>ClockA,
            CD=>scuba_vlo, Q=>addr010_ff);

    FF_7: FD1P3DX
        -- synopsys translate_off
        generic map (GSR=> "ENABLED")
        -- synopsys translate_on
        port map (D=>AddressA(11), SP=>wren0_inv_g, CK=>ClockA,
            CD=>scuba_vlo, Q=>addr011_ff);

    FF_6: FD1P3DX
        -- synopsys translate_off
        generic map (GSR=> "ENABLED")
        -- synopsys translate_on
        port map (D=>AddressA(12), SP=>wren0_inv_g, CK=>ClockA,
            CD=>scuba_vlo, Q=>addr012_ff);

    FF_5: FD1P3DX
        -- synopsys translate_off
        generic map (GSR=> "ENABLED")
        -- synopsys translate_on
        port map (D=>AddressB(10), SP=>wren1_inv_g, CK=>ClockB,
            CD=>scuba_vlo, Q=>addr110_ff);

    FF_4: FD1P3DX
        -- synopsys translate_off
        generic map (GSR=> "ENABLED")
        -- synopsys translate_on
        port map (D=>AddressB(11), SP=>wren1_inv_g, CK=>ClockB,
            CD=>scuba_vlo, Q=>addr111_ff);

    FF_3: FD1P3DX
        -- synopsys translate_off
        generic map (GSR=> "ENABLED")
        -- synopsys translate_on
        port map (D=>AddressB(12), SP=>wren1_inv_g, CK=>ClockB,
            CD=>scuba_vlo, Q=>addr112_ff);

    FF_2: FD1P3DX
        -- synopsys translate_off
        generic map (GSR=> "ENABLED")
        -- synopsys translate_on
        port map (D=>addr110_ff, SP=>ClockEnB, CK=>ClockB, CD=>scuba_vlo,
            Q=>addr110_ff2);

    FF_1: FD1P3DX
        -- synopsys translate_off
        generic map (GSR=> "ENABLED")
        -- synopsys translate_on
        port map (D=>addr111_ff, SP=>ClockEnB, CK=>ClockB, CD=>scuba_vlo,
            Q=>addr111_ff2);

    FF_0: FD1P3DX
        -- synopsys translate_off
        generic map (GSR=> "ENABLED")
        -- synopsys translate_on
        port map (D=>addr112_ff, SP=>ClockEnB, CK=>ClockB, CD=>scuba_vlo,
            Q=>addr112_ff2);

    mux_31: MUX81
        port map (D0=>mdout0_0_0, D1=>mdout0_1_0, D2=>mdout0_2_0,
            D3=>mdout0_3_0, D4=>mdout0_4_0, D5=>mdout0_5_0,
            D6=>scuba_vlo, D7=>scuba_vlo, SD1=>addr010_ff,
            SD2=>addr011_ff, SD3=>addr012_ff, Z=>QA(0));

    mux_30: MUX81
        port map (D0=>mdout0_0_1, D1=>mdout0_1_1, D2=>mdout0_2_1,
            D3=>mdout0_3_1, D4=>mdout0_4_1, D5=>mdout0_5_1,
            D6=>scuba_vlo, D7=>scuba_vlo, SD1=>addr010_ff,
            SD2=>addr011_ff, SD3=>addr012_ff, Z=>QA(1));

    mux_29: MUX81
        port map (D0=>mdout0_0_2, D1=>mdout0_1_2, D2=>mdout0_2_2,
            D3=>mdout0_3_2, D4=>mdout0_4_2, D5=>mdout0_5_2,
            D6=>scuba_vlo, D7=>scuba_vlo, SD1=>addr010_ff,
            SD2=>addr011_ff, SD3=>addr012_ff, Z=>QA(2));

    mux_28: MUX81
        port map (D0=>mdout0_0_3, D1=>mdout0_1_3, D2=>mdout0_2_3,
            D3=>mdout0_3_3, D4=>mdout0_4_3, D5=>mdout0_5_3,
            D6=>scuba_vlo, D7=>scuba_vlo, SD1=>addr010_ff,
            SD2=>addr011_ff, SD3=>addr012_ff, Z=>QA(3));

    mux_27: MUX81
        port map (D0=>mdout0_0_4, D1=>mdout0_1_4, D2=>mdout0_2_4,
            D3=>mdout0_3_4, D4=>mdout0_4_4, D5=>mdout0_5_4,
            D6=>scuba_vlo, D7=>scuba_vlo, SD1=>addr010_ff,
            SD2=>addr011_ff, SD3=>addr012_ff, Z=>QA(4));

    mux_26: MUX81
        port map (D0=>mdout0_0_5, D1=>mdout0_1_5, D2=>mdout0_2_5,
            D3=>mdout0_3_5, D4=>mdout0_4_5, D5=>mdout0_5_5,
            D6=>scuba_vlo, D7=>scuba_vlo, SD1=>addr010_ff,
            SD2=>addr011_ff, SD3=>addr012_ff, Z=>QA(5));

    mux_25: MUX81
        port map (D0=>mdout0_0_6, D1=>mdout0_1_6, D2=>mdout0_2_6,
            D3=>mdout0_3_6, D4=>mdout0_4_6, D5=>mdout0_5_6,
            D6=>scuba_vlo, D7=>scuba_vlo, SD1=>addr010_ff,
            SD2=>addr011_ff, SD3=>addr012_ff, Z=>QA(6));

    mux_24: MUX81
        port map (D0=>mdout0_0_7, D1=>mdout0_1_7, D2=>mdout0_2_7,
            D3=>mdout0_3_7, D4=>mdout0_4_7, D5=>mdout0_5_7,
            D6=>scuba_vlo, D7=>scuba_vlo, SD1=>addr010_ff,
            SD2=>addr011_ff, SD3=>addr012_ff, Z=>QA(7));

    mux_23: MUX81
        port map (D0=>mdout0_0_9, D1=>mdout0_1_9, D2=>mdout0_2_9,
            D3=>mdout0_3_9, D4=>mdout0_4_9, D5=>mdout0_5_9,
            D6=>scuba_vlo, D7=>scuba_vlo, SD1=>addr010_ff,
            SD2=>addr011_ff, SD3=>addr012_ff, Z=>QA(8));

    mux_22: MUX81
        port map (D0=>mdout0_0_10, D1=>mdout0_1_10, D2=>mdout0_2_10,
            D3=>mdout0_3_10, D4=>mdout0_4_10, D5=>mdout0_5_10,
            D6=>scuba_vlo, D7=>scuba_vlo, SD1=>addr010_ff,
            SD2=>addr011_ff, SD3=>addr012_ff, Z=>QA(9));

    mux_21: MUX81
        port map (D0=>mdout0_0_11, D1=>mdout0_1_11, D2=>mdout0_2_11,
            D3=>mdout0_3_11, D4=>mdout0_4_11, D5=>mdout0_5_11,
            D6=>scuba_vlo, D7=>scuba_vlo, SD1=>addr010_ff,
            SD2=>addr011_ff, SD3=>addr012_ff, Z=>QA(10));

    mux_20: MUX81
        port map (D0=>mdout0_0_12, D1=>mdout0_1_12, D2=>mdout0_2_12,
            D3=>mdout0_3_12, D4=>mdout0_4_12, D5=>mdout0_5_12,
            D6=>scuba_vlo, D7=>scuba_vlo, SD1=>addr010_ff,
            SD2=>addr011_ff, SD3=>addr012_ff, Z=>QA(11));

    mux_19: MUX81
        port map (D0=>mdout0_0_13, D1=>mdout0_1_13, D2=>mdout0_2_13,
            D3=>mdout0_3_13, D4=>mdout0_4_13, D5=>mdout0_5_13,
            D6=>scuba_vlo, D7=>scuba_vlo, SD1=>addr010_ff,
            SD2=>addr011_ff, SD3=>addr012_ff, Z=>QA(12));

    mux_18: MUX81
        port map (D0=>mdout0_0_14, D1=>mdout0_1_14, D2=>mdout0_2_14,
            D3=>mdout0_3_14, D4=>mdout0_4_14, D5=>mdout0_5_14,
            D6=>scuba_vlo, D7=>scuba_vlo, SD1=>addr010_ff,
            SD2=>addr011_ff, SD3=>addr012_ff, Z=>QA(13));

    mux_17: MUX81
        port map (D0=>mdout0_0_15, D1=>mdout0_1_15, D2=>mdout0_2_15,
            D3=>mdout0_3_15, D4=>mdout0_4_15, D5=>mdout0_5_15,
            D6=>scuba_vlo, D7=>scuba_vlo, SD1=>addr010_ff,
            SD2=>addr011_ff, SD3=>addr012_ff, Z=>QA(14));

    mux_16: MUX81
        port map (D0=>mdout0_0_16, D1=>mdout0_1_16, D2=>mdout0_2_16,
            D3=>mdout0_3_16, D4=>mdout0_4_16, D5=>mdout0_5_16,
            D6=>scuba_vlo, D7=>scuba_vlo, SD1=>addr010_ff,
            SD2=>addr011_ff, SD3=>addr012_ff, Z=>QA(15));

    mux_15: MUX81
        port map (D0=>mdout1_0_0, D1=>mdout1_1_0, D2=>mdout1_2_0,
            D3=>mdout1_3_0, D4=>mdout1_4_0, D5=>mdout1_5_0,
            D6=>scuba_vlo, D7=>scuba_vlo, SD1=>addr110_ff2,
            SD2=>addr111_ff2, SD3=>addr112_ff2, Z=>QB(0));

    mux_14: MUX81
        port map (D0=>mdout1_0_1, D1=>mdout1_1_1, D2=>mdout1_2_1,
            D3=>mdout1_3_1, D4=>mdout1_4_1, D5=>mdout1_5_1,
            D6=>scuba_vlo, D7=>scuba_vlo, SD1=>addr110_ff2,
            SD2=>addr111_ff2, SD3=>addr112_ff2, Z=>QB(1));

    mux_13: MUX81
        port map (D0=>mdout1_0_2, D1=>mdout1_1_2, D2=>mdout1_2_2,
            D3=>mdout1_3_2, D4=>mdout1_4_2, D5=>mdout1_5_2,
            D6=>scuba_vlo, D7=>scuba_vlo, SD1=>addr110_ff2,
            SD2=>addr111_ff2, SD3=>addr112_ff2, Z=>QB(2));

    mux_12: MUX81
        port map (D0=>mdout1_0_3, D1=>mdout1_1_3, D2=>mdout1_2_3,
            D3=>mdout1_3_3, D4=>mdout1_4_3, D5=>mdout1_5_3,
            D6=>scuba_vlo, D7=>scuba_vlo, SD1=>addr110_ff2,
            SD2=>addr111_ff2, SD3=>addr112_ff2, Z=>QB(3));

    mux_11: MUX81
        port map (D0=>mdout1_0_4, D1=>mdout1_1_4, D2=>mdout1_2_4,
            D3=>mdout1_3_4, D4=>mdout1_4_4, D5=>mdout1_5_4,
            D6=>scuba_vlo, D7=>scuba_vlo, SD1=>addr110_ff2,
            SD2=>addr111_ff2, SD3=>addr112_ff2, Z=>QB(4));

    mux_10: MUX81
        port map (D0=>mdout1_0_5, D1=>mdout1_1_5, D2=>mdout1_2_5,
            D3=>mdout1_3_5, D4=>mdout1_4_5, D5=>mdout1_5_5,
            D6=>scuba_vlo, D7=>scuba_vlo, SD1=>addr110_ff2,
            SD2=>addr111_ff2, SD3=>addr112_ff2, Z=>QB(5));

    mux_9: MUX81
        port map (D0=>mdout1_0_6, D1=>mdout1_1_6, D2=>mdout1_2_6,
            D3=>mdout1_3_6, D4=>mdout1_4_6, D5=>mdout1_5_6,
            D6=>scuba_vlo, D7=>scuba_vlo, SD1=>addr110_ff2,
            SD2=>addr111_ff2, SD3=>addr112_ff2, Z=>QB(6));

    mux_8: MUX81
        port map (D0=>mdout1_0_7, D1=>mdout1_1_7, D2=>mdout1_2_7,
            D3=>mdout1_3_7, D4=>mdout1_4_7, D5=>mdout1_5_7,
            D6=>scuba_vlo, D7=>scuba_vlo, SD1=>addr110_ff2,
            SD2=>addr111_ff2, SD3=>addr112_ff2, Z=>QB(7));

    mux_7: MUX81
        port map (D0=>mdout1_0_9, D1=>mdout1_1_9, D2=>mdout1_2_9,
            D3=>mdout1_3_9, D4=>mdout1_4_9, D5=>mdout1_5_9,
            D6=>scuba_vlo, D7=>scuba_vlo, SD1=>addr110_ff2,
            SD2=>addr111_ff2, SD3=>addr112_ff2, Z=>QB(8));

    mux_6: MUX81
        port map (D0=>mdout1_0_10, D1=>mdout1_1_10, D2=>mdout1_2_10,
            D3=>mdout1_3_10, D4=>mdout1_4_10, D5=>mdout1_5_10,
            D6=>scuba_vlo, D7=>scuba_vlo, SD1=>addr110_ff2,
            SD2=>addr111_ff2, SD3=>addr112_ff2, Z=>QB(9));

    mux_5: MUX81
        port map (D0=>mdout1_0_11, D1=>mdout1_1_11, D2=>mdout1_2_11,
            D3=>mdout1_3_11, D4=>mdout1_4_11, D5=>mdout1_5_11,
            D6=>scuba_vlo, D7=>scuba_vlo, SD1=>addr110_ff2,
            SD2=>addr111_ff2, SD3=>addr112_ff2, Z=>QB(10));

    mux_4: MUX81
        port map (D0=>mdout1_0_12, D1=>mdout1_1_12, D2=>mdout1_2_12,
            D3=>mdout1_3_12, D4=>mdout1_4_12, D5=>mdout1_5_12,
            D6=>scuba_vlo, D7=>scuba_vlo, SD1=>addr110_ff2,
            SD2=>addr111_ff2, SD3=>addr112_ff2, Z=>QB(11));

    mux_3: MUX81
        port map (D0=>mdout1_0_13, D1=>mdout1_1_13, D2=>mdout1_2_13,
            D3=>mdout1_3_13, D4=>mdout1_4_13, D5=>mdout1_5_13,
            D6=>scuba_vlo, D7=>scuba_vlo, SD1=>addr110_ff2,
            SD2=>addr111_ff2, SD3=>addr112_ff2, Z=>QB(12));

    mux_2: MUX81
        port map (D0=>mdout1_0_14, D1=>mdout1_1_14, D2=>mdout1_2_14,
            D3=>mdout1_3_14, D4=>mdout1_4_14, D5=>mdout1_5_14,
            D6=>scuba_vlo, D7=>scuba_vlo, SD1=>addr110_ff2,
            SD2=>addr111_ff2, SD3=>addr112_ff2, Z=>QB(13));

    mux_1: MUX81
        port map (D0=>mdout1_0_15, D1=>mdout1_1_15, D2=>mdout1_2_15,
            D3=>mdout1_3_15, D4=>mdout1_4_15, D5=>mdout1_5_15,
            D6=>scuba_vlo, D7=>scuba_vlo, SD1=>addr110_ff2,
            SD2=>addr111_ff2, SD3=>addr112_ff2, Z=>QB(14));

    scuba_vlo_inst: VLO
        port map (Z=>scuba_vlo);

    mux_0: MUX81
        port map (D0=>mdout1_0_16, D1=>mdout1_1_16, D2=>mdout1_2_16,
            D3=>mdout1_3_16, D4=>mdout1_4_16, D5=>mdout1_5_16,
            D6=>scuba_vlo, D7=>scuba_vlo, SD1=>addr110_ff2,
            SD2=>addr111_ff2, SD3=>addr112_ff2, Z=>QB(15));

end Structure;

-- synopsys translate_off
library xp2;
configuration Structure_CON of byte_cache_16 is
    for Structure
        for all:AND2 use entity xp2.AND2(V); end for;
        for all:FD1P3DX use entity xp2.FD1P3DX(V); end for;
        for all:INV use entity xp2.INV(V); end for;
        for all:MUX81 use entity xp2.MUX81(V); end for;
        for all:VHI use entity xp2.VHI(V); end for;
        for all:VLO use entity xp2.VLO(V); end for;
        for all:DP16KB use entity xp2.DP16KB(V); end for;
    end for;
end Structure_CON;

-- synopsys translate_on