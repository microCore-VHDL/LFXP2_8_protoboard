-- ---------------------------------------------------------------------
-- @file : debugger.vhd
-- ---------------------------------------------------------------------
--
-- Last change: KS 15.12.2020 17:07:54
-- Project : microCore
-- Language : VHDL-2008
-- Last check in : $Rev: 612 $ $Date:: 2020-12-16 #$
-- @copyright (c): Klaus Schleisiek, All Rights Reserved.
--
-- Do not use this file except in compliance with the License. You may
-- obtain a copy of the License at http://www.microcore.org/License/.
-- Software distributed under the License is distributed on an "AS IS"
-- basis, WITHOUT WARRANTY OF ANY KIND, either express or implied.
-- See the License for the specific language governing rights and
-- limitations under the License.
--
-- @brief: The debugger connects to the host via an RS232 interface
--         and allows interactive control while microCore is running.
--         The debugger does not use the processor, it is a specific
--         set of state machines.
--
-- Version Author   Date       Changes
--           ks    8-Jun-2020  initial version
-- ---------------------------------------------------------------------
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_signed.ALL;
USE work.functions_pkg.ALL;
USE work.architecture_pkg.ALL;

ENTITY debugger IS PORT (
   uBus           : IN  uBus_port;
   deb_reset      : OUT STD_LOGIC;    -- reset generated by debugger
   deb_pause      : OUT STD_LOGIC;
   deb_prequest   : OUT STD_LOGIC;    -- request program memory write cycle
   deb_penable    : IN  STD_LOGIC;    -- execute program memory write
   deb_drequest   : OUT STD_LOGIC;    -- request data memory for a read/write cycle
   deb_denable    : IN  STD_LOGIC;    -- execute data memory read/write
   umbilical      : OUT progmem_port; -- interface to the program memory
   debugmem       : OUT datamem_port; -- interface to the data memory
   debugmem_rdata : IN  data_bus;
-- umbilical uart
   rxd            : IN  STD_LOGIC;
   break          : OUT STD_LOGIC;
   txd            : OUT STD_LOGIC
); END debugger;

ARCHITECTURE rtl OF debugger IS

CONSTANT addr_width   : NATURAL := max(data_addr_width, prog_addr_width);

ALIAS  reset       : STD_LOGIC IS uBus.reset;
ALIAS  clk         : STD_LOGIC IS uBus.clk;
ALIAS  clk_en      : STD_LOGIC IS uBus.clk_en;
ALIAS  wdata       : data_bus  IS uBus.wdata;
SIGNAL progload    : STD_LOGIC;

COMPONENT uart GENERIC (
   rate       : NATURAL;
   depth      : NATURAL;
   ramstyle   : STRING
); PORT (
   uBus       : IN  uBus_port;
   pause      : OUT STD_LOGIC; -- uart pause
   rx_full    : OUT STD_LOGIC; -- rx data buffer full
   rx_read    : IN  STD_LOGIC; -- read rx data buffer
   rx_data    : OUT byte;      -- rx data buffer
   rx_break   : OUT STD_LOGIC; -- break detected
   rx_ovrn    : OUT STD_LOGIC; -- rx overrun, queue = full+1
   tx_empty   : OUT STD_LOGIC; -- data buffer empty
   tx_write   : IN  STD_LOGIC; -- write into data buffer
   tx_data    : IN  byte;      -- output data
   tx_busy    : OUT STD_LOGIC; -- tx uart still busy
-- UART I/O
   dtr        : IN  STD_LOGIC;
   rxd        : IN  STD_LOGIC;
   txd        : OUT STD_LOGIC
); END COMPONENT uart;

SIGNAL rx_full     : STD_LOGIC;  -- uart buffer full
SIGNAL rx_read     : STD_LOGIC;  -- read uart buffer
SIGNAL rx_data     : byte;       -- uart input buffer
SIGNAL tx_empty    : STD_LOGIC;  -- uart buffer empty
SIGNAL tx_write    : STD_LOGIC;  -- write byte
SIGNAL tx_data     : byte;       -- uart output buffer
SIGNAL uart_break  : STD_LOGIC;  -- break from uart
SIGNAL host_break  : STD_LOGIC;  -- break via umbilical

-- umbilical
CONSTANT all_nibbles : STD_LOGIC_VECTOR(log2(octetts)-1 DOWNTO 0) := to_vec(octetts-1, log2(octetts));

-- umbilical uart input
TYPE in_states     IS (idle, getaddr, getlength, loading, rx_debug, full, ack, uploading, downloading);

SIGNAL in_state    : in_states;
SIGNAL in_ctr      : STD_LOGIC_VECTOR(log2(octetts)-1 DOWNTO 0); -- #nibbles to receive from host
SIGNAL in_reg      : STD_LOGIC_VECTOR(octetts*8-1 DOWNTO 0);
SIGNAL in_rd       : STD_LOGIC;  -- target reads in_reg
SIGNAL upload      : STD_LOGIC;
SIGNAL download    : STD_LOGIC;
SIGNAL addr_ptr    : STD_LOGIC_VECTOR(addr_width-1 DOWNTO 0);
SIGNAL addr_ctr    : STD_LOGIC_VECTOR(addr_width-1 DOWNTO 0);

-- umbilical uart output
TYPE out_states    IS (start, idle, mark, tx_debug, wait_ack, readmem, downloading);

SIGNAL out_state   : out_states;
SIGNAL out_ctr     : STD_LOGIC_VECTOR(log2(octetts)-1 DOWNTO 0); -- #nibbles to receive from host
SIGNAL out_wr      : STD_LOGIC;  -- target writes out_reg
SIGNAL out_reg     : STD_LOGIC_VECTOR(octetts*8-1 DOWNTO 0);
SIGNAL send_ack    : STD_LOGIC;

-- memory control
SIGNAL dread       : STD_LOGIC;
SIGNAL write       : STD_LOGIC;  -- write signal for umbilical

-- pragma translate_off
SIGNAL in_read     : STD_LOGIC;
SIGNAL out_written : STD_LOGIC;
-- pragma translate_on

BEGIN

break        <= host_break OR uart_break;
deb_prequest <= write AND progload;

-- pragma translate_off
in_read     <= '0' WHEN  in_state /= full                       ELSE in_rd;  -- for simulation only
out_written <= '0' WHEN  out_state /= idle OR in_state /= idle  ELSE out_wr; -- for simulation only
-- pragma translate_on

umbilical.enable <= deb_penable;
umbilical.write  <= write;
umbilical.read   <= '0';
umbilical.addr   <= addr_ptr(prog_addr_width-1 DOWNTO 0);
umbilical.wdata  <= rx_data;

debugmem.enable  <= deb_denable WHEN  with_up_download  ELSE '0';
debugmem.write   <= write;
debugmem.addr    <= addr_ptr(data_addr_width-1 DOWNTO 0);
debugmem.wdata   <= in_reg(data_width-1 DOWNTO 0);

in_rd  <= '1' WHEN  uReg_read (uBus, DEBUG_REG)  ELSE '0';
out_wr <= '1' WHEN  uReg_write(uBus, DEBUG_REG)  ELSE '0';

deb_pause <= '1' WHEN  (in_rd  = '1' AND  in_state /= full) OR
                       (out_wr = '1' AND (in_state /= idle OR out_state /= idle))
                 ELSE '0';

-- ---------------------------------------------------------------------
-- loading the program memory
-- and listening to the host
-- ---------------------------------------------------------------------

tx_data <= mark_ack   WHEN  send_ack = '1'     ELSE
           mark_debug WHEN  out_state = mark   ELSE
           mark_nack  WHEN  out_state = start  ELSE
           out_reg(out_reg'high DOWNTO out_reg'high-7);

umbilical_proc: PROCESS(clk, reset)

   PROCEDURE tx_ack IS
   BEGIN
      IF  out_state = idle AND tx_empty = '1' AND tx_write = '0'  THEN
         send_ack <= '1';
         tx_write <= '1';
      END IF;
   END tx_ack;

   PROCEDURE tx_start IS
   BEGIN
      IF  tx_empty = '1' AND tx_write = '0'  THEN
         tx_write <= '1';
      END IF;
   END tx_start;

BEGIN
   IF  reset = '1' AND async_reset  THEN
         out_ctr <= all_nibbles;
       out_state <= start;
        in_state <= idle;
        progload <= '0';
        send_ack <= '0';
          upload <= '0';
        download <= '0';
      host_break <= '0';
           write <= '0';
       deb_reset <= '0';
    deb_drequest <= '0';
   ELSIF  rising_edge(clk)  THEN
      IF  clk_en = '1'  THEN
         tx_write <= '0';
         dread <= '0';

         IF  deb_penable = '1'  THEN
            addr_ptr <= addr_ptr + 1;
            addr_ctr <= addr_ctr - 1;
         END IF;

         IF  deb_denable = '1'  THEN
            dread <= '1';
            write <= '0';
            deb_drequest <= '0';
            addr_ptr <= addr_ptr + 1;
            addr_ctr <= addr_ctr - 1;
         END IF;

-- ---------------------------------------------------------------------
-- umbilical input
-- ---------------------------------------------------------------------

         CASE in_state IS

         WHEN idle      => in_ctr <= all_nibbles;
                           progload <= '0';
                           upload <= '0';
                           IF  rx_full = '1' AND download = '0'  THEN
                              CASE rx_data IS
                              WHEN mark_start    => in_state <= getaddr;
                                                    progload <= '1';
                              WHEN mark_reset    => deb_reset <= '1';
                                                    in_state <= getaddr;
                                                    progload <= '1';
                              WHEN mark_debug    => in_state <= rx_debug;
                              WHEN mark_upload   => IF  with_up_download  THEN
                                                       in_state <= getaddr;
                                                       upload <= '1';
                                                    END IF;
                              WHEN mark_download => IF  with_up_download  THEN
                                                       in_state <= getaddr;
                                                       download <= '1';
                                                    END IF;
                              WHEN mark_break    => host_break <= '1';
                              WHEN mark_nbreak   => host_break <= '0';
                              WHEN OTHERS        => NULL;
                              END CASE;
                           END IF;

         WHEN getaddr   => IF  rx_full = '1'  THEN
                              in_reg <= in_reg(in_reg'high-8 DOWNTO 0) & rx_data;
                              in_ctr <= in_ctr - 1;
                              IF  in_ctr = 0  THEN
                                 in_ctr <= all_nibbles;
                                 addr_ptr <= in_reg(addr_width-9 DOWNTO 0) & rx_data;
                                 in_state <= getlength;
                              END IF;
                           END IF;

         WHEN getlength => IF  rx_full = '1'  THEN
                              in_reg <= in_reg(in_reg'high-8 DOWNTO 0) & rx_data;
                              in_ctr <= in_ctr - 1;
                              IF  in_ctr = 0  THEN
                                 in_ctr <= all_nibbles;
                                 addr_ctr <= in_reg(addr_width-9 DOWNTO 0) & rx_data;
                                 in_state <= loading;
                                 IF  upload = '1' AND with_up_download  THEN
                                    in_state <= uploading;
                                 END IF;
                                 IF  download = '1' AND with_up_download  THEN
                                    in_state <= downloading;
                                 END IF;
                              END IF;
                           END IF;

         WHEN loading   => IF  addr_ctr = 0  THEN
                              tx_ack;
                              IF  send_ack = '1'  THEN
                                 send_ack <= '0';
                                 in_state <= idle;
                                 deb_reset <= '0';
                              END IF;
                           ELSIF  rx_full = '1'  THEN
                              write <= '1';
                           ELSIF  deb_penable = '1'  THEN
                              write <= '0';
                           END IF;

         WHEN rx_debug  => IF  rx_full = '1'  THEN
                              in_reg <= in_reg(in_reg'high-8 DOWNTO 0) & rx_data;
                              in_ctr <= in_ctr - 1;
                              IF  in_ctr = 0  THEN
                                 in_ctr <= all_nibbles;
                                 in_state <= full;
                              END IF;
                           END IF;

         WHEN full      => IF  in_rd = '1'  THEN
                              in_state <= ack;
                           END IF;

         WHEN ack       => tx_ack;
                           IF  send_ack = '1'  THEN
                              send_ack <= '0';
                              in_state <= idle;
                           END IF;

         WHEN uploading => IF  with_up_download  THEN
                              IF  addr_ctr = 0  THEN
                                 tx_ack;
                                 IF  send_ack = '1'  THEN
                                    send_ack <= '0';
                                    in_state <= idle;
                                 END IF;
                              ELSIF  rx_full = '1'  THEN
                                 in_reg <= in_reg(in_reg'high-8 DOWNTO 0) & rx_data;
                                 IF  in_ctr = 0  THEN
                                    in_ctr <= all_nibbles;
                                    deb_drequest <= '1';
                                    write <= '1';
                                 ELSE
                                    in_ctr <= in_ctr - 1;
                                 END IF;
                              END IF;
                           END IF;

         WHEN downloading => IF  with_up_download  THEN
                              IF  out_state = idle  THEN
                                 deb_drequest <= '1';
                                 out_state <= readmem;
                                 in_state <= idle;
                              END IF;
                           END IF;

         WHEN OTHERS    => in_state <= idle;

         END CASE;

-- ---------------------------------------------------------------------
-- umbilical output
-- ---------------------------------------------------------------------

         CASE out_state IS

         WHEN start     => tx_start;
                           IF  tx_write = '1'  THEN
                              IF  out_ctr = 0  THEN
                                 out_state <= idle;
                              ELSE
                                 out_ctr <= out_ctr - 1;
                              END IF;
                           END IF;

         WHEN idle      => out_ctr <= all_nibbles;
                           IF  out_wr = '1' AND in_state = idle AND send_ack = '0'  THEN   -- send a new word
                              out_reg <= to_vec(0, out_reg'length - data_width) & wdata;
                              out_state <= mark;
                           END IF;

         WHEN mark      => tx_start;
                           IF  tx_write = '1'  THEN
                              out_state <= tx_debug;
                           END IF;

         WHEN tx_debug  => tx_start;
                           IF  tx_write = '1'  THEN
                              IF  out_ctr = 0  THEN
                                 out_state <= wait_ack;
                              ELSE
                                 out_reg <= out_reg(out_reg'high-8 DOWNTO 0) & "00000000";
                                 out_ctr <= out_ctr - 1;
                              END IF;
                           END IF;

         WHEN wait_ack  => IF  rx_full = '1' AND rx_data = mark_ack  THEN
                              out_state <= idle;
                              download <= '0';
                           END IF;

         WHEN readmem   => IF  with_up_download  THEN
                              IF  dread = '1'  THEN
                                 out_reg <= to_vec(0, out_reg'length - data_width) & debugmem_rdata;
                                 out_ctr <= all_nibbles;
                                 out_state <= downloading;
                              END IF;
                           END IF;

         WHEN downloading => IF  with_up_download  THEN
                              tx_start;
                              IF  tx_write = '1'  THEN
                                 IF  out_ctr /= 0  THEN
                                    out_reg <= out_reg(out_reg'high-8 DOWNTO 0) & "00000000";
                                    out_ctr <= out_ctr - 1;
                                 ELSIF  addr_ctr /= 0  THEN
                                    deb_drequest <= '1';
                                    out_state <= readmem;
                                 ELSE -- addr_ctr = 0
                                    out_state <= wait_ack;
                                 END IF;
                              END IF;
                           END IF;

         WHEN OTHERS    => out_state <= idle;

         END CASE;

      END IF; -- clk_en = '1'

      IF  reset = '1' AND NOT async_reset  THEN
           out_ctr <= all_nibbles;
         out_state <= start;
          in_state <= idle;
          progload <= '0';
          send_ack <= '0';
            upload <= '0';
          download <= '0';
        host_break <= '0';
             write <= '0';
         deb_reset <= '0';
      deb_drequest <= '0';
      END IF;

   END IF;
END PROCESS umbilical_proc;

-- ---------------------------------------------------------------------
-- umbilical uart
-- ---------------------------------------------------------------------

rx_read <= rx_full AND clk_en;

debug_uart: uart
GENERIC MAP (umbilical_rate, 4, "registers") PORT MAP (
   uBus       => uBus,
   pause      => OPEN,
   rx_full    => rx_full,    -- rx data buffer full
   rx_read    => rx_read,    -- read rx data buffer
   rx_data    => rx_data,    -- rx data buffer
   rx_break   => uart_break, -- break detected
   rx_ovrn    => OPEN,
   tx_empty   => tx_empty,   -- data buffer empty
   tx_write   => tx_write,   -- write into data buffer
   tx_data    => tx_data,    -- output data
   tx_busy    => OPEN,
-- UART I/O
   dtr        => '1',
   rxd        => rxd,
   txd        => txd
);

END rtl;